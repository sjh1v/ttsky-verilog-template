magic
tech sky130A
magscale 1 2
timestamp 1765482302
<< checkpaint >>
rect -1260 8332 31260 31260
rect -1486 -172 31260 8332
rect -1260 -1260 31260 -172
<< viali >>
rect 1501 27557 1535 27591
rect 7297 27557 7331 27591
rect 25237 27489 25271 27523
rect 16221 27421 16255 27455
rect 25513 27421 25547 27455
rect 1777 27353 1811 27387
rect 7573 27353 7607 27387
rect 16405 27285 16439 27319
rect 28273 25245 28307 25279
rect 28549 25245 28583 25279
rect 1409 18717 1443 18751
rect 1685 18717 1719 18751
rect 16681 13277 16715 13311
rect 16037 13141 16071 13175
rect 15853 12937 15887 12971
rect 15945 12937 15979 12971
rect 17049 12869 17083 12903
rect 16497 12801 16531 12835
rect 17141 12801 17175 12835
rect 17509 12801 17543 12835
rect 18429 12801 18463 12835
rect 19257 12801 19291 12835
rect 16129 12733 16163 12767
rect 17325 12733 17359 12767
rect 18061 12733 18095 12767
rect 18337 12733 18371 12767
rect 19165 12733 19199 12767
rect 16681 12665 16715 12699
rect 18797 12665 18831 12699
rect 18889 12665 18923 12699
rect 15485 12597 15519 12631
rect 16313 12597 16347 12631
rect 18153 12325 18187 12359
rect 15945 12257 15979 12291
rect 17877 12257 17911 12291
rect 15117 12189 15151 12223
rect 15669 12189 15703 12223
rect 17785 12189 17819 12223
rect 14933 12053 14967 12087
rect 17417 12053 17451 12087
rect 17601 11849 17635 11883
rect 14657 11781 14691 11815
rect 17693 11713 17727 11747
rect 18061 11713 18095 11747
rect 18981 11713 19015 11747
rect 19625 11713 19659 11747
rect 14381 11645 14415 11679
rect 17785 11645 17819 11679
rect 18613 11645 18647 11679
rect 18889 11645 18923 11679
rect 19809 11645 19843 11679
rect 20177 11645 20211 11679
rect 16129 11577 16163 11611
rect 19349 11577 19383 11611
rect 17233 11509 17267 11543
rect 19441 11509 19475 11543
rect 21603 11509 21637 11543
rect 13829 11305 13863 11339
rect 19257 11305 19291 11339
rect 21005 11305 21039 11339
rect 17969 11237 18003 11271
rect 13461 11169 13495 11203
rect 14473 11169 14507 11203
rect 19809 11169 19843 11203
rect 13553 11101 13587 11135
rect 14197 11101 14231 11135
rect 16221 11101 16255 11135
rect 18981 11101 19015 11135
rect 19625 11101 19659 11135
rect 20729 11101 20763 11135
rect 22753 11101 22787 11135
rect 16497 11033 16531 11067
rect 19717 11033 19751 11067
rect 20085 11033 20119 11067
rect 22477 11033 22511 11067
rect 15945 10965 15979 10999
rect 18429 10965 18463 10999
rect 14565 10761 14599 10795
rect 14933 10761 14967 10795
rect 15025 10761 15059 10795
rect 17325 10761 17359 10795
rect 17877 10761 17911 10795
rect 18337 10761 18371 10795
rect 20453 10761 20487 10795
rect 21465 10761 21499 10795
rect 24685 10693 24719 10727
rect 15209 10625 15243 10659
rect 16865 10625 16899 10659
rect 17509 10625 17543 10659
rect 17969 10625 18003 10659
rect 18613 10625 18647 10659
rect 21281 10625 21315 10659
rect 21925 10625 21959 10659
rect 22201 10625 22235 10659
rect 22293 10625 22327 10659
rect 14381 10557 14415 10591
rect 14473 10557 14507 10591
rect 15301 10557 15335 10591
rect 15945 10557 15979 10591
rect 16773 10557 16807 10591
rect 17785 10557 17819 10591
rect 18705 10557 18739 10591
rect 18981 10557 19015 10591
rect 22661 10557 22695 10591
rect 22937 10557 22971 10591
rect 17233 10489 17267 10523
rect 21925 10489 21959 10523
rect 22477 10489 22511 10523
rect 18429 10421 18463 10455
rect 14105 10081 14139 10115
rect 16957 10081 16991 10115
rect 17233 10081 17267 10115
rect 18705 10081 18739 10115
rect 20545 10081 20579 10115
rect 21557 10081 21591 10115
rect 22201 10081 22235 10115
rect 16589 10013 16623 10047
rect 20085 10013 20119 10047
rect 21097 10013 21131 10047
rect 21189 10013 21223 10047
rect 21833 10013 21867 10047
rect 22017 10013 22051 10047
rect 14381 9945 14415 9979
rect 20177 9945 20211 9979
rect 20269 9945 20303 9979
rect 20407 9945 20441 9979
rect 21465 9945 21499 9979
rect 22477 9945 22511 9979
rect 24225 9945 24259 9979
rect 15853 9877 15887 9911
rect 15945 9877 15979 9911
rect 19901 9877 19935 9911
rect 20913 9877 20947 9911
rect 21649 9877 21683 9911
rect 14933 9673 14967 9707
rect 19625 9673 19659 9707
rect 22201 9673 22235 9707
rect 23029 9673 23063 9707
rect 21097 9605 21131 9639
rect 14381 9537 14415 9571
rect 14473 9537 14507 9571
rect 15117 9537 15151 9571
rect 15485 9537 15519 9571
rect 17417 9537 17451 9571
rect 18429 9537 18463 9571
rect 19165 9537 19199 9571
rect 19809 9537 19843 9571
rect 20821 9537 20855 9571
rect 21005 9537 21039 9571
rect 21189 9537 21223 9571
rect 21925 9537 21959 9571
rect 22569 9537 22603 9571
rect 23213 9537 23247 9571
rect 23305 9537 23339 9571
rect 23581 9537 23615 9571
rect 14197 9469 14231 9503
rect 15577 9469 15611 9503
rect 15853 9469 15887 9503
rect 17555 9469 17589 9503
rect 17693 9469 17727 9503
rect 18613 9469 18647 9503
rect 19901 9469 19935 9503
rect 19993 9469 20027 9503
rect 20085 9469 20119 9503
rect 20545 9469 20579 9503
rect 20637 9469 20671 9503
rect 20729 9469 20763 9503
rect 22017 9469 22051 9503
rect 22661 9469 22695 9503
rect 22753 9469 22787 9503
rect 23673 9469 23707 9503
rect 14841 9401 14875 9435
rect 17969 9401 18003 9435
rect 20361 9401 20395 9435
rect 16773 9333 16807 9367
rect 19257 9333 19291 9367
rect 20269 9333 20303 9367
rect 18337 9129 18371 9163
rect 20453 9129 20487 9163
rect 20913 9129 20947 9163
rect 21097 9129 21131 9163
rect 22109 9129 22143 9163
rect 22293 9129 22327 9163
rect 14381 9061 14415 9095
rect 23029 9061 23063 9095
rect 15025 8993 15059 9027
rect 15945 8993 15979 9027
rect 16497 8993 16531 9027
rect 17141 8993 17175 9027
rect 17417 8993 17451 9027
rect 17534 8993 17568 9027
rect 17693 8993 17727 9027
rect 20729 8993 20763 9027
rect 21649 8993 21683 9027
rect 1409 8925 1443 8959
rect 14289 8925 14323 8959
rect 16037 8925 16071 8959
rect 16681 8925 16715 8959
rect 18429 8925 18463 8959
rect 18613 8925 18647 8959
rect 19349 8925 19383 8959
rect 20085 8925 20119 8959
rect 21005 8925 21039 8959
rect 21465 8925 21499 8959
rect 22385 8925 22419 8959
rect 23121 8925 23155 8959
rect 23305 8925 23339 8959
rect 23581 8925 23615 8959
rect 24685 8925 24719 8959
rect 14749 8857 14783 8891
rect 20269 8857 20303 8891
rect 21925 8857 21959 8891
rect 22141 8857 22175 8891
rect 22870 8857 22904 8891
rect 1593 8789 1627 8823
rect 14105 8789 14139 8823
rect 14841 8789 14875 8823
rect 15301 8789 15335 8823
rect 16221 8789 16255 8823
rect 18429 8789 18463 8823
rect 19993 8789 20027 8823
rect 20729 8789 20763 8823
rect 21557 8789 21591 8823
rect 22661 8789 22695 8823
rect 22753 8789 22787 8823
rect 23765 8789 23799 8823
rect 24501 8789 24535 8823
rect 15669 8585 15703 8619
rect 16681 8585 16715 8619
rect 18245 8585 18279 8619
rect 21373 8585 21407 8619
rect 22845 8585 22879 8619
rect 23213 8585 23247 8619
rect 14197 8517 14231 8551
rect 16313 8517 16347 8551
rect 17049 8517 17083 8551
rect 22937 8517 22971 8551
rect 23029 8517 23063 8551
rect 23581 8517 23615 8551
rect 13921 8449 13955 8483
rect 15945 8449 15979 8483
rect 17141 8449 17175 8483
rect 17509 8449 17543 8483
rect 19993 8449 20027 8483
rect 20269 8449 20303 8483
rect 20361 8449 20395 8483
rect 20637 8449 20671 8483
rect 20821 8449 20855 8483
rect 20913 8449 20947 8483
rect 21281 8449 21315 8483
rect 21649 8449 21683 8483
rect 21833 8449 21867 8483
rect 22477 8449 22511 8483
rect 22661 8449 22695 8483
rect 17325 8381 17359 8415
rect 18061 8381 18095 8415
rect 19717 8381 19751 8415
rect 20085 8381 20119 8415
rect 20545 8381 20579 8415
rect 21189 8381 21223 8415
rect 23305 8381 23339 8415
rect 21925 8313 21959 8347
rect 25053 8313 25087 8347
rect 15945 8041 15979 8075
rect 19257 8041 19291 8075
rect 20545 8041 20579 8075
rect 23765 8041 23799 8075
rect 23949 8041 23983 8075
rect 24501 8041 24535 8075
rect 19901 7973 19935 8007
rect 18153 7905 18187 7939
rect 18981 7905 19015 7939
rect 19993 7905 20027 7939
rect 24133 7905 24167 7939
rect 17417 7837 17451 7871
rect 17693 7837 17727 7871
rect 17785 7837 17819 7871
rect 17877 7837 17911 7871
rect 18705 7837 18739 7871
rect 19533 7837 19567 7871
rect 19625 7837 19659 7871
rect 21833 7837 21867 7871
rect 23949 7837 23983 7871
rect 24409 7837 24443 7871
rect 24685 7837 24719 7871
rect 24961 7837 24995 7871
rect 18015 7769 18049 7803
rect 18797 7769 18831 7803
rect 21925 7769 21959 7803
rect 24225 7769 24259 7803
rect 17509 7701 17543 7735
rect 18337 7701 18371 7735
rect 19717 7701 19751 7735
rect 23213 7701 23247 7735
rect 24869 7701 24903 7735
rect 25145 7701 25179 7735
rect 14749 7497 14783 7531
rect 17601 7497 17635 7531
rect 18337 7497 18371 7531
rect 20545 7497 20579 7531
rect 20713 7497 20747 7531
rect 21097 7497 21131 7531
rect 22477 7497 22511 7531
rect 16221 7429 16255 7463
rect 17233 7429 17267 7463
rect 17417 7429 17451 7463
rect 20453 7429 20487 7463
rect 20913 7429 20947 7463
rect 21465 7429 21499 7463
rect 17693 7361 17727 7395
rect 21189 7361 21223 7395
rect 21649 7361 21683 7395
rect 21833 7361 21867 7395
rect 21925 7361 21959 7395
rect 22109 7361 22143 7395
rect 22201 7361 22235 7395
rect 22293 7361 22327 7395
rect 16497 7293 16531 7327
rect 18429 7293 18463 7327
rect 18705 7293 18739 7327
rect 22569 7293 22603 7327
rect 22753 7293 22787 7327
rect 22845 7293 22879 7327
rect 22937 7293 22971 7327
rect 23029 7293 23063 7327
rect 23397 7293 23431 7327
rect 23673 7293 23707 7327
rect 20729 7157 20763 7191
rect 21281 7157 21315 7191
rect 25145 7157 25179 7191
rect 16668 6953 16702 6987
rect 18153 6953 18187 6987
rect 18705 6953 18739 6987
rect 21575 6953 21609 6987
rect 23305 6953 23339 6987
rect 23397 6953 23431 6987
rect 25329 6953 25363 6987
rect 21833 6817 21867 6851
rect 24961 6817 24995 6851
rect 16405 6749 16439 6783
rect 18521 6749 18555 6783
rect 18981 6749 19015 6783
rect 21925 6749 21959 6783
rect 22569 6749 22603 6783
rect 23029 6749 23063 6783
rect 23121 6749 23155 6783
rect 23581 6749 23615 6783
rect 23765 6749 23799 6783
rect 23949 6749 23983 6783
rect 24409 6749 24443 6783
rect 25421 6749 25455 6783
rect 25697 6749 25731 6783
rect 23673 6681 23707 6715
rect 18797 6613 18831 6647
rect 20085 6613 20119 6647
rect 22661 6613 22695 6647
rect 25145 6613 25179 6647
rect 20361 6409 20395 6443
rect 22661 6409 22695 6443
rect 23213 6409 23247 6443
rect 23857 6409 23891 6443
rect 19993 6341 20027 6375
rect 22845 6341 22879 6375
rect 23121 6341 23155 6375
rect 20545 6273 20579 6307
rect 21005 6273 21039 6307
rect 21189 6273 21223 6307
rect 22293 6273 22327 6307
rect 22385 6273 22419 6307
rect 23029 6273 23063 6307
rect 23581 6273 23615 6307
rect 23765 6273 23799 6307
rect 24041 6273 24075 6307
rect 28273 6273 28307 6307
rect 16681 6205 16715 6239
rect 16957 6205 16991 6239
rect 18429 6205 18463 6239
rect 20269 6205 20303 6239
rect 23397 6205 23431 6239
rect 24225 6205 24259 6239
rect 24501 6205 24535 6239
rect 25973 6205 26007 6239
rect 26709 6205 26743 6239
rect 28549 6205 28583 6239
rect 21189 6137 21223 6171
rect 26157 6137 26191 6171
rect 18521 6069 18555 6103
rect 22477 6069 22511 6103
rect 19073 5865 19107 5899
rect 23489 5865 23523 5899
rect 24409 5865 24443 5899
rect 17601 5729 17635 5763
rect 18153 5729 18187 5763
rect 18613 5729 18647 5763
rect 18705 5729 18739 5763
rect 19257 5729 19291 5763
rect 19809 5729 19843 5763
rect 20453 5729 20487 5763
rect 22017 5729 22051 5763
rect 23305 5729 23339 5763
rect 23949 5729 23983 5763
rect 24685 5729 24719 5763
rect 25053 5729 25087 5763
rect 18429 5661 18463 5695
rect 18889 5661 18923 5695
rect 20177 5661 20211 5695
rect 22202 5639 22236 5673
rect 22385 5661 22419 5695
rect 22661 5661 22695 5695
rect 22753 5661 22787 5695
rect 23673 5661 23707 5695
rect 23765 5661 23799 5695
rect 23857 5661 23891 5695
rect 24593 5661 24627 5695
rect 25145 5661 25179 5695
rect 25421 5661 25455 5695
rect 25605 5661 25639 5695
rect 17417 5593 17451 5627
rect 22293 5593 22327 5627
rect 22503 5593 22537 5627
rect 16129 5525 16163 5559
rect 18245 5525 18279 5559
rect 21925 5525 21959 5559
rect 25329 5525 25363 5559
rect 19717 5321 19751 5355
rect 20269 5321 20303 5355
rect 22477 5321 22511 5355
rect 22937 5321 22971 5355
rect 23397 5321 23431 5355
rect 16957 5253 16991 5287
rect 19809 5253 19843 5287
rect 25237 5253 25271 5287
rect 19257 5185 19291 5219
rect 19533 5185 19567 5219
rect 20085 5185 20119 5219
rect 20545 5185 20579 5219
rect 21373 5185 21407 5219
rect 21833 5185 21867 5219
rect 22477 5185 22511 5219
rect 22569 5185 22603 5219
rect 22753 5185 22787 5219
rect 23121 5185 23155 5219
rect 23581 5185 23615 5219
rect 23673 5185 23707 5219
rect 23765 5185 23799 5219
rect 23857 5185 23891 5219
rect 24133 5185 24167 5219
rect 24317 5185 24351 5219
rect 24409 5185 24443 5219
rect 24501 5185 24535 5219
rect 24777 5185 24811 5219
rect 24961 5185 24995 5219
rect 16681 5117 16715 5151
rect 18429 5117 18463 5151
rect 19073 5117 19107 5151
rect 19349 5117 19383 5151
rect 19993 5117 20027 5151
rect 20729 5117 20763 5151
rect 20821 5117 20855 5151
rect 23305 5117 23339 5151
rect 25881 5117 25915 5151
rect 22017 5049 22051 5083
rect 24777 5049 24811 5083
rect 18521 4981 18555 5015
rect 19349 4981 19383 5015
rect 19809 4981 19843 5015
rect 20361 4981 20395 5015
rect 24685 4981 24719 5015
rect 17785 4777 17819 4811
rect 18705 4777 18739 4811
rect 21005 4777 21039 4811
rect 26157 4777 26191 4811
rect 18981 4709 19015 4743
rect 15853 4641 15887 4675
rect 17601 4641 17635 4675
rect 18153 4641 18187 4675
rect 24409 4641 24443 4675
rect 24685 4641 24719 4675
rect 17969 4573 18003 4607
rect 18797 4573 18831 4607
rect 19257 4573 19291 4607
rect 21281 4573 21315 4607
rect 21465 4573 21499 4607
rect 21557 4573 21591 4607
rect 21741 4573 21775 4607
rect 22109 4573 22143 4607
rect 22753 4573 22787 4607
rect 23673 4573 23707 4607
rect 16129 4505 16163 4539
rect 19533 4505 19567 4539
rect 22845 4505 22879 4539
rect 23029 4505 23063 4539
rect 21097 4437 21131 4471
rect 21925 4437 21959 4471
rect 22661 4437 22695 4471
rect 22937 4437 22971 4471
rect 23581 4437 23615 4471
rect 16313 4233 16347 4267
rect 19441 4233 19475 4267
rect 21557 4233 21591 4267
rect 22569 4233 22603 4267
rect 23949 4233 23983 4267
rect 24961 4233 24995 4267
rect 22109 4165 22143 4199
rect 22201 4165 22235 4199
rect 22339 4165 22373 4199
rect 22753 4165 22787 4199
rect 16497 4097 16531 4131
rect 17417 4097 17451 4131
rect 17877 4097 17911 4131
rect 18981 4097 19015 4131
rect 19165 4097 19199 4131
rect 19349 4097 19383 4131
rect 19625 4097 19659 4131
rect 22017 4097 22051 4131
rect 22477 4097 22511 4131
rect 22845 4097 22879 4131
rect 22937 4097 22971 4131
rect 23213 4097 23247 4131
rect 23489 4097 23523 4131
rect 23946 4097 23980 4131
rect 17601 4029 17635 4063
rect 17693 4029 17727 4063
rect 18889 4029 18923 4063
rect 19809 4029 19843 4063
rect 20085 4029 20119 4063
rect 21833 4029 21867 4063
rect 23305 4029 23339 4063
rect 24317 4029 24351 4063
rect 24409 4029 24443 4063
rect 25605 4029 25639 4063
rect 18245 3961 18279 3995
rect 23121 3961 23155 3995
rect 17233 3893 17267 3927
rect 18061 3893 18095 3927
rect 23397 3893 23431 3927
rect 23673 3893 23707 3927
rect 23765 3893 23799 3927
rect 18337 3689 18371 3723
rect 23121 3689 23155 3723
rect 26157 3689 26191 3723
rect 23581 3621 23615 3655
rect 16589 3553 16623 3587
rect 19901 3553 19935 3587
rect 20177 3553 20211 3587
rect 22569 3553 22603 3587
rect 24409 3553 24443 3587
rect 24685 3553 24719 3587
rect 18889 3485 18923 3519
rect 20269 3485 20303 3519
rect 20361 3485 20395 3519
rect 20821 3485 20855 3519
rect 22845 3485 22879 3519
rect 23213 3485 23247 3519
rect 23305 3485 23339 3519
rect 23397 3485 23431 3519
rect 23581 3485 23615 3519
rect 16865 3417 16899 3451
rect 18521 3417 18555 3451
rect 19257 3349 19291 3383
rect 20729 3349 20763 3383
rect 22661 3349 22695 3383
rect 17233 3145 17267 3179
rect 19625 3145 19659 3179
rect 18153 3077 18187 3111
rect 17417 3009 17451 3043
rect 17877 3009 17911 3043
rect 19717 3009 19751 3043
rect 21833 3009 21867 3043
rect 19993 2941 20027 2975
rect 22109 2941 22143 2975
rect 23581 2941 23615 2975
rect 24225 2941 24259 2975
rect 21465 2873 21499 2907
rect 23673 2805 23707 2839
rect 18153 2601 18187 2635
rect 20269 2601 20303 2635
rect 21189 2601 21223 2635
rect 22017 2601 22051 2635
rect 22753 2601 22787 2635
rect 19717 2533 19751 2567
rect 23029 2533 23063 2567
rect 1685 2465 1719 2499
rect 19349 2465 19383 2499
rect 22201 2465 22235 2499
rect 22661 2465 22695 2499
rect 1409 2397 1443 2431
rect 9137 2397 9171 2431
rect 18337 2397 18371 2431
rect 19533 2397 19567 2431
rect 20453 2397 20487 2431
rect 21281 2397 21315 2431
rect 22293 2397 22327 2431
rect 23029 2397 23063 2431
rect 23213 2397 23247 2431
rect 27353 2397 27387 2431
rect 9321 2261 9355 2295
rect 27169 2261 27203 2295
<< metal1 >>
rect 1104 27770 28888 27792
rect 1104 27718 4423 27770
rect 4475 27718 4487 27770
rect 4539 27718 4551 27770
rect 4603 27718 4615 27770
rect 4667 27718 4679 27770
rect 4731 27718 11369 27770
rect 11421 27718 11433 27770
rect 11485 27718 11497 27770
rect 11549 27718 11561 27770
rect 11613 27718 11625 27770
rect 11677 27718 18315 27770
rect 18367 27718 18379 27770
rect 18431 27718 18443 27770
rect 18495 27718 18507 27770
rect 18559 27718 18571 27770
rect 18623 27718 25261 27770
rect 25313 27718 25325 27770
rect 25377 27718 25389 27770
rect 25441 27718 25453 27770
rect 25505 27718 25517 27770
rect 25569 27718 28888 27770
rect 1104 27696 28888 27718
rect 16040 27628 16252 27656
rect 1486 27548 1492 27600
rect 1544 27548 1550 27600
rect 7190 27548 7196 27600
rect 7248 27588 7254 27600
rect 7285 27591 7343 27597
rect 7285 27588 7297 27591
rect 7248 27560 7297 27588
rect 7248 27548 7254 27560
rect 7285 27557 7297 27560
rect 7331 27557 7343 27591
rect 16040 27588 16068 27628
rect 7285 27551 7343 27557
rect 7484 27560 16068 27588
rect 1765 27387 1823 27393
rect 1765 27353 1777 27387
rect 1811 27384 1823 27387
rect 7484 27384 7512 27560
rect 16114 27548 16120 27600
rect 16172 27548 16178 27600
rect 16224 27588 16252 27628
rect 21634 27588 21640 27600
rect 16224 27560 21640 27588
rect 21634 27548 21640 27560
rect 21692 27548 21698 27600
rect 16132 27452 16160 27548
rect 25130 27480 25136 27532
rect 25188 27520 25194 27532
rect 25225 27523 25283 27529
rect 25225 27520 25237 27523
rect 25188 27492 25237 27520
rect 25188 27480 25194 27492
rect 25225 27489 25237 27492
rect 25271 27489 25283 27523
rect 25225 27483 25283 27489
rect 16209 27455 16267 27461
rect 16209 27452 16221 27455
rect 16132 27424 16221 27452
rect 16209 27421 16221 27424
rect 16255 27421 16267 27455
rect 16209 27415 16267 27421
rect 17586 27412 17592 27464
rect 17644 27452 17650 27464
rect 25501 27455 25559 27461
rect 25501 27452 25513 27455
rect 17644 27424 25513 27452
rect 17644 27412 17650 27424
rect 25501 27421 25513 27424
rect 25547 27421 25559 27455
rect 25501 27415 25559 27421
rect 7561 27387 7619 27393
rect 7561 27384 7573 27387
rect 1811 27356 6914 27384
rect 7484 27356 7573 27384
rect 1811 27353 1823 27356
rect 1765 27347 1823 27353
rect 6886 27316 6914 27356
rect 7561 27353 7573 27356
rect 7607 27353 7619 27387
rect 20990 27384 20996 27396
rect 7561 27347 7619 27353
rect 7668 27356 20996 27384
rect 7668 27316 7696 27356
rect 20990 27344 20996 27356
rect 21048 27344 21054 27396
rect 6886 27288 7696 27316
rect 15838 27276 15844 27328
rect 15896 27316 15902 27328
rect 16393 27319 16451 27325
rect 16393 27316 16405 27319
rect 15896 27288 16405 27316
rect 15896 27276 15902 27288
rect 16393 27285 16405 27288
rect 16439 27285 16451 27319
rect 16393 27279 16451 27285
rect 1104 27226 28888 27248
rect 1104 27174 5083 27226
rect 5135 27174 5147 27226
rect 5199 27174 5211 27226
rect 5263 27174 5275 27226
rect 5327 27174 5339 27226
rect 5391 27174 12029 27226
rect 12081 27174 12093 27226
rect 12145 27174 12157 27226
rect 12209 27174 12221 27226
rect 12273 27174 12285 27226
rect 12337 27174 18975 27226
rect 19027 27174 19039 27226
rect 19091 27174 19103 27226
rect 19155 27174 19167 27226
rect 19219 27174 19231 27226
rect 19283 27174 25921 27226
rect 25973 27174 25985 27226
rect 26037 27174 26049 27226
rect 26101 27174 26113 27226
rect 26165 27174 26177 27226
rect 26229 27174 28888 27226
rect 1104 27152 28888 27174
rect 1104 26682 28888 26704
rect 1104 26630 4423 26682
rect 4475 26630 4487 26682
rect 4539 26630 4551 26682
rect 4603 26630 4615 26682
rect 4667 26630 4679 26682
rect 4731 26630 11369 26682
rect 11421 26630 11433 26682
rect 11485 26630 11497 26682
rect 11549 26630 11561 26682
rect 11613 26630 11625 26682
rect 11677 26630 18315 26682
rect 18367 26630 18379 26682
rect 18431 26630 18443 26682
rect 18495 26630 18507 26682
rect 18559 26630 18571 26682
rect 18623 26630 25261 26682
rect 25313 26630 25325 26682
rect 25377 26630 25389 26682
rect 25441 26630 25453 26682
rect 25505 26630 25517 26682
rect 25569 26630 28888 26682
rect 1104 26608 28888 26630
rect 1104 26138 28888 26160
rect 1104 26086 5083 26138
rect 5135 26086 5147 26138
rect 5199 26086 5211 26138
rect 5263 26086 5275 26138
rect 5327 26086 5339 26138
rect 5391 26086 12029 26138
rect 12081 26086 12093 26138
rect 12145 26086 12157 26138
rect 12209 26086 12221 26138
rect 12273 26086 12285 26138
rect 12337 26086 18975 26138
rect 19027 26086 19039 26138
rect 19091 26086 19103 26138
rect 19155 26086 19167 26138
rect 19219 26086 19231 26138
rect 19283 26086 25921 26138
rect 25973 26086 25985 26138
rect 26037 26086 26049 26138
rect 26101 26086 26113 26138
rect 26165 26086 26177 26138
rect 26229 26086 28888 26138
rect 1104 26064 28888 26086
rect 1104 25594 28888 25616
rect 1104 25542 4423 25594
rect 4475 25542 4487 25594
rect 4539 25542 4551 25594
rect 4603 25542 4615 25594
rect 4667 25542 4679 25594
rect 4731 25542 11369 25594
rect 11421 25542 11433 25594
rect 11485 25542 11497 25594
rect 11549 25542 11561 25594
rect 11613 25542 11625 25594
rect 11677 25542 18315 25594
rect 18367 25542 18379 25594
rect 18431 25542 18443 25594
rect 18495 25542 18507 25594
rect 18559 25542 18571 25594
rect 18623 25542 25261 25594
rect 25313 25542 25325 25594
rect 25377 25542 25389 25594
rect 25441 25542 25453 25594
rect 25505 25542 25517 25594
rect 25569 25542 28888 25594
rect 1104 25520 28888 25542
rect 28258 25236 28264 25288
rect 28316 25236 28322 25288
rect 28534 25236 28540 25288
rect 28592 25236 28598 25288
rect 1104 25050 28888 25072
rect 1104 24998 5083 25050
rect 5135 24998 5147 25050
rect 5199 24998 5211 25050
rect 5263 24998 5275 25050
rect 5327 24998 5339 25050
rect 5391 24998 12029 25050
rect 12081 24998 12093 25050
rect 12145 24998 12157 25050
rect 12209 24998 12221 25050
rect 12273 24998 12285 25050
rect 12337 24998 18975 25050
rect 19027 24998 19039 25050
rect 19091 24998 19103 25050
rect 19155 24998 19167 25050
rect 19219 24998 19231 25050
rect 19283 24998 25921 25050
rect 25973 24998 25985 25050
rect 26037 24998 26049 25050
rect 26101 24998 26113 25050
rect 26165 24998 26177 25050
rect 26229 24998 28888 25050
rect 1104 24976 28888 24998
rect 1104 24506 28888 24528
rect 1104 24454 4423 24506
rect 4475 24454 4487 24506
rect 4539 24454 4551 24506
rect 4603 24454 4615 24506
rect 4667 24454 4679 24506
rect 4731 24454 11369 24506
rect 11421 24454 11433 24506
rect 11485 24454 11497 24506
rect 11549 24454 11561 24506
rect 11613 24454 11625 24506
rect 11677 24454 18315 24506
rect 18367 24454 18379 24506
rect 18431 24454 18443 24506
rect 18495 24454 18507 24506
rect 18559 24454 18571 24506
rect 18623 24454 25261 24506
rect 25313 24454 25325 24506
rect 25377 24454 25389 24506
rect 25441 24454 25453 24506
rect 25505 24454 25517 24506
rect 25569 24454 28888 24506
rect 1104 24432 28888 24454
rect 1104 23962 28888 23984
rect 1104 23910 5083 23962
rect 5135 23910 5147 23962
rect 5199 23910 5211 23962
rect 5263 23910 5275 23962
rect 5327 23910 5339 23962
rect 5391 23910 12029 23962
rect 12081 23910 12093 23962
rect 12145 23910 12157 23962
rect 12209 23910 12221 23962
rect 12273 23910 12285 23962
rect 12337 23910 18975 23962
rect 19027 23910 19039 23962
rect 19091 23910 19103 23962
rect 19155 23910 19167 23962
rect 19219 23910 19231 23962
rect 19283 23910 25921 23962
rect 25973 23910 25985 23962
rect 26037 23910 26049 23962
rect 26101 23910 26113 23962
rect 26165 23910 26177 23962
rect 26229 23910 28888 23962
rect 1104 23888 28888 23910
rect 1104 23418 28888 23440
rect 1104 23366 4423 23418
rect 4475 23366 4487 23418
rect 4539 23366 4551 23418
rect 4603 23366 4615 23418
rect 4667 23366 4679 23418
rect 4731 23366 11369 23418
rect 11421 23366 11433 23418
rect 11485 23366 11497 23418
rect 11549 23366 11561 23418
rect 11613 23366 11625 23418
rect 11677 23366 18315 23418
rect 18367 23366 18379 23418
rect 18431 23366 18443 23418
rect 18495 23366 18507 23418
rect 18559 23366 18571 23418
rect 18623 23366 25261 23418
rect 25313 23366 25325 23418
rect 25377 23366 25389 23418
rect 25441 23366 25453 23418
rect 25505 23366 25517 23418
rect 25569 23366 28888 23418
rect 1104 23344 28888 23366
rect 1104 22874 28888 22896
rect 1104 22822 5083 22874
rect 5135 22822 5147 22874
rect 5199 22822 5211 22874
rect 5263 22822 5275 22874
rect 5327 22822 5339 22874
rect 5391 22822 12029 22874
rect 12081 22822 12093 22874
rect 12145 22822 12157 22874
rect 12209 22822 12221 22874
rect 12273 22822 12285 22874
rect 12337 22822 18975 22874
rect 19027 22822 19039 22874
rect 19091 22822 19103 22874
rect 19155 22822 19167 22874
rect 19219 22822 19231 22874
rect 19283 22822 25921 22874
rect 25973 22822 25985 22874
rect 26037 22822 26049 22874
rect 26101 22822 26113 22874
rect 26165 22822 26177 22874
rect 26229 22822 28888 22874
rect 1104 22800 28888 22822
rect 1104 22330 28888 22352
rect 1104 22278 4423 22330
rect 4475 22278 4487 22330
rect 4539 22278 4551 22330
rect 4603 22278 4615 22330
rect 4667 22278 4679 22330
rect 4731 22278 11369 22330
rect 11421 22278 11433 22330
rect 11485 22278 11497 22330
rect 11549 22278 11561 22330
rect 11613 22278 11625 22330
rect 11677 22278 18315 22330
rect 18367 22278 18379 22330
rect 18431 22278 18443 22330
rect 18495 22278 18507 22330
rect 18559 22278 18571 22330
rect 18623 22278 25261 22330
rect 25313 22278 25325 22330
rect 25377 22278 25389 22330
rect 25441 22278 25453 22330
rect 25505 22278 25517 22330
rect 25569 22278 28888 22330
rect 1104 22256 28888 22278
rect 1104 21786 28888 21808
rect 1104 21734 5083 21786
rect 5135 21734 5147 21786
rect 5199 21734 5211 21786
rect 5263 21734 5275 21786
rect 5327 21734 5339 21786
rect 5391 21734 12029 21786
rect 12081 21734 12093 21786
rect 12145 21734 12157 21786
rect 12209 21734 12221 21786
rect 12273 21734 12285 21786
rect 12337 21734 18975 21786
rect 19027 21734 19039 21786
rect 19091 21734 19103 21786
rect 19155 21734 19167 21786
rect 19219 21734 19231 21786
rect 19283 21734 25921 21786
rect 25973 21734 25985 21786
rect 26037 21734 26049 21786
rect 26101 21734 26113 21786
rect 26165 21734 26177 21786
rect 26229 21734 28888 21786
rect 1104 21712 28888 21734
rect 1104 21242 28888 21264
rect 1104 21190 4423 21242
rect 4475 21190 4487 21242
rect 4539 21190 4551 21242
rect 4603 21190 4615 21242
rect 4667 21190 4679 21242
rect 4731 21190 11369 21242
rect 11421 21190 11433 21242
rect 11485 21190 11497 21242
rect 11549 21190 11561 21242
rect 11613 21190 11625 21242
rect 11677 21190 18315 21242
rect 18367 21190 18379 21242
rect 18431 21190 18443 21242
rect 18495 21190 18507 21242
rect 18559 21190 18571 21242
rect 18623 21190 25261 21242
rect 25313 21190 25325 21242
rect 25377 21190 25389 21242
rect 25441 21190 25453 21242
rect 25505 21190 25517 21242
rect 25569 21190 28888 21242
rect 1104 21168 28888 21190
rect 1104 20698 28888 20720
rect 1104 20646 5083 20698
rect 5135 20646 5147 20698
rect 5199 20646 5211 20698
rect 5263 20646 5275 20698
rect 5327 20646 5339 20698
rect 5391 20646 12029 20698
rect 12081 20646 12093 20698
rect 12145 20646 12157 20698
rect 12209 20646 12221 20698
rect 12273 20646 12285 20698
rect 12337 20646 18975 20698
rect 19027 20646 19039 20698
rect 19091 20646 19103 20698
rect 19155 20646 19167 20698
rect 19219 20646 19231 20698
rect 19283 20646 25921 20698
rect 25973 20646 25985 20698
rect 26037 20646 26049 20698
rect 26101 20646 26113 20698
rect 26165 20646 26177 20698
rect 26229 20646 28888 20698
rect 1104 20624 28888 20646
rect 1104 20154 28888 20176
rect 1104 20102 4423 20154
rect 4475 20102 4487 20154
rect 4539 20102 4551 20154
rect 4603 20102 4615 20154
rect 4667 20102 4679 20154
rect 4731 20102 11369 20154
rect 11421 20102 11433 20154
rect 11485 20102 11497 20154
rect 11549 20102 11561 20154
rect 11613 20102 11625 20154
rect 11677 20102 18315 20154
rect 18367 20102 18379 20154
rect 18431 20102 18443 20154
rect 18495 20102 18507 20154
rect 18559 20102 18571 20154
rect 18623 20102 25261 20154
rect 25313 20102 25325 20154
rect 25377 20102 25389 20154
rect 25441 20102 25453 20154
rect 25505 20102 25517 20154
rect 25569 20102 28888 20154
rect 1104 20080 28888 20102
rect 1104 19610 28888 19632
rect 1104 19558 5083 19610
rect 5135 19558 5147 19610
rect 5199 19558 5211 19610
rect 5263 19558 5275 19610
rect 5327 19558 5339 19610
rect 5391 19558 12029 19610
rect 12081 19558 12093 19610
rect 12145 19558 12157 19610
rect 12209 19558 12221 19610
rect 12273 19558 12285 19610
rect 12337 19558 18975 19610
rect 19027 19558 19039 19610
rect 19091 19558 19103 19610
rect 19155 19558 19167 19610
rect 19219 19558 19231 19610
rect 19283 19558 25921 19610
rect 25973 19558 25985 19610
rect 26037 19558 26049 19610
rect 26101 19558 26113 19610
rect 26165 19558 26177 19610
rect 26229 19558 28888 19610
rect 1104 19536 28888 19558
rect 1104 19066 28888 19088
rect 1104 19014 4423 19066
rect 4475 19014 4487 19066
rect 4539 19014 4551 19066
rect 4603 19014 4615 19066
rect 4667 19014 4679 19066
rect 4731 19014 11369 19066
rect 11421 19014 11433 19066
rect 11485 19014 11497 19066
rect 11549 19014 11561 19066
rect 11613 19014 11625 19066
rect 11677 19014 18315 19066
rect 18367 19014 18379 19066
rect 18431 19014 18443 19066
rect 18495 19014 18507 19066
rect 18559 19014 18571 19066
rect 18623 19014 25261 19066
rect 25313 19014 25325 19066
rect 25377 19014 25389 19066
rect 25441 19014 25453 19066
rect 25505 19014 25517 19066
rect 25569 19014 28888 19066
rect 1104 18992 28888 19014
rect 934 18708 940 18760
rect 992 18748 998 18760
rect 1397 18751 1455 18757
rect 1397 18748 1409 18751
rect 992 18720 1409 18748
rect 992 18708 998 18720
rect 1397 18717 1409 18720
rect 1443 18717 1455 18751
rect 1397 18711 1455 18717
rect 1673 18751 1731 18757
rect 1673 18717 1685 18751
rect 1719 18748 1731 18751
rect 13446 18748 13452 18760
rect 1719 18720 13452 18748
rect 1719 18717 1731 18720
rect 1673 18711 1731 18717
rect 13446 18708 13452 18720
rect 13504 18708 13510 18760
rect 1104 18522 28888 18544
rect 1104 18470 5083 18522
rect 5135 18470 5147 18522
rect 5199 18470 5211 18522
rect 5263 18470 5275 18522
rect 5327 18470 5339 18522
rect 5391 18470 12029 18522
rect 12081 18470 12093 18522
rect 12145 18470 12157 18522
rect 12209 18470 12221 18522
rect 12273 18470 12285 18522
rect 12337 18470 18975 18522
rect 19027 18470 19039 18522
rect 19091 18470 19103 18522
rect 19155 18470 19167 18522
rect 19219 18470 19231 18522
rect 19283 18470 25921 18522
rect 25973 18470 25985 18522
rect 26037 18470 26049 18522
rect 26101 18470 26113 18522
rect 26165 18470 26177 18522
rect 26229 18470 28888 18522
rect 1104 18448 28888 18470
rect 1104 17978 28888 18000
rect 1104 17926 4423 17978
rect 4475 17926 4487 17978
rect 4539 17926 4551 17978
rect 4603 17926 4615 17978
rect 4667 17926 4679 17978
rect 4731 17926 11369 17978
rect 11421 17926 11433 17978
rect 11485 17926 11497 17978
rect 11549 17926 11561 17978
rect 11613 17926 11625 17978
rect 11677 17926 18315 17978
rect 18367 17926 18379 17978
rect 18431 17926 18443 17978
rect 18495 17926 18507 17978
rect 18559 17926 18571 17978
rect 18623 17926 25261 17978
rect 25313 17926 25325 17978
rect 25377 17926 25389 17978
rect 25441 17926 25453 17978
rect 25505 17926 25517 17978
rect 25569 17926 28888 17978
rect 1104 17904 28888 17926
rect 1104 17434 28888 17456
rect 1104 17382 5083 17434
rect 5135 17382 5147 17434
rect 5199 17382 5211 17434
rect 5263 17382 5275 17434
rect 5327 17382 5339 17434
rect 5391 17382 12029 17434
rect 12081 17382 12093 17434
rect 12145 17382 12157 17434
rect 12209 17382 12221 17434
rect 12273 17382 12285 17434
rect 12337 17382 18975 17434
rect 19027 17382 19039 17434
rect 19091 17382 19103 17434
rect 19155 17382 19167 17434
rect 19219 17382 19231 17434
rect 19283 17382 25921 17434
rect 25973 17382 25985 17434
rect 26037 17382 26049 17434
rect 26101 17382 26113 17434
rect 26165 17382 26177 17434
rect 26229 17382 28888 17434
rect 1104 17360 28888 17382
rect 1104 16890 28888 16912
rect 1104 16838 4423 16890
rect 4475 16838 4487 16890
rect 4539 16838 4551 16890
rect 4603 16838 4615 16890
rect 4667 16838 4679 16890
rect 4731 16838 11369 16890
rect 11421 16838 11433 16890
rect 11485 16838 11497 16890
rect 11549 16838 11561 16890
rect 11613 16838 11625 16890
rect 11677 16838 18315 16890
rect 18367 16838 18379 16890
rect 18431 16838 18443 16890
rect 18495 16838 18507 16890
rect 18559 16838 18571 16890
rect 18623 16838 25261 16890
rect 25313 16838 25325 16890
rect 25377 16838 25389 16890
rect 25441 16838 25453 16890
rect 25505 16838 25517 16890
rect 25569 16838 28888 16890
rect 1104 16816 28888 16838
rect 1104 16346 28888 16368
rect 1104 16294 5083 16346
rect 5135 16294 5147 16346
rect 5199 16294 5211 16346
rect 5263 16294 5275 16346
rect 5327 16294 5339 16346
rect 5391 16294 12029 16346
rect 12081 16294 12093 16346
rect 12145 16294 12157 16346
rect 12209 16294 12221 16346
rect 12273 16294 12285 16346
rect 12337 16294 18975 16346
rect 19027 16294 19039 16346
rect 19091 16294 19103 16346
rect 19155 16294 19167 16346
rect 19219 16294 19231 16346
rect 19283 16294 25921 16346
rect 25973 16294 25985 16346
rect 26037 16294 26049 16346
rect 26101 16294 26113 16346
rect 26165 16294 26177 16346
rect 26229 16294 28888 16346
rect 1104 16272 28888 16294
rect 1104 15802 28888 15824
rect 1104 15750 4423 15802
rect 4475 15750 4487 15802
rect 4539 15750 4551 15802
rect 4603 15750 4615 15802
rect 4667 15750 4679 15802
rect 4731 15750 11369 15802
rect 11421 15750 11433 15802
rect 11485 15750 11497 15802
rect 11549 15750 11561 15802
rect 11613 15750 11625 15802
rect 11677 15750 18315 15802
rect 18367 15750 18379 15802
rect 18431 15750 18443 15802
rect 18495 15750 18507 15802
rect 18559 15750 18571 15802
rect 18623 15750 25261 15802
rect 25313 15750 25325 15802
rect 25377 15750 25389 15802
rect 25441 15750 25453 15802
rect 25505 15750 25517 15802
rect 25569 15750 28888 15802
rect 1104 15728 28888 15750
rect 1104 15258 28888 15280
rect 1104 15206 5083 15258
rect 5135 15206 5147 15258
rect 5199 15206 5211 15258
rect 5263 15206 5275 15258
rect 5327 15206 5339 15258
rect 5391 15206 12029 15258
rect 12081 15206 12093 15258
rect 12145 15206 12157 15258
rect 12209 15206 12221 15258
rect 12273 15206 12285 15258
rect 12337 15206 18975 15258
rect 19027 15206 19039 15258
rect 19091 15206 19103 15258
rect 19155 15206 19167 15258
rect 19219 15206 19231 15258
rect 19283 15206 25921 15258
rect 25973 15206 25985 15258
rect 26037 15206 26049 15258
rect 26101 15206 26113 15258
rect 26165 15206 26177 15258
rect 26229 15206 28888 15258
rect 1104 15184 28888 15206
rect 1104 14714 28888 14736
rect 1104 14662 4423 14714
rect 4475 14662 4487 14714
rect 4539 14662 4551 14714
rect 4603 14662 4615 14714
rect 4667 14662 4679 14714
rect 4731 14662 11369 14714
rect 11421 14662 11433 14714
rect 11485 14662 11497 14714
rect 11549 14662 11561 14714
rect 11613 14662 11625 14714
rect 11677 14662 18315 14714
rect 18367 14662 18379 14714
rect 18431 14662 18443 14714
rect 18495 14662 18507 14714
rect 18559 14662 18571 14714
rect 18623 14662 25261 14714
rect 25313 14662 25325 14714
rect 25377 14662 25389 14714
rect 25441 14662 25453 14714
rect 25505 14662 25517 14714
rect 25569 14662 28888 14714
rect 1104 14640 28888 14662
rect 1104 14170 28888 14192
rect 1104 14118 5083 14170
rect 5135 14118 5147 14170
rect 5199 14118 5211 14170
rect 5263 14118 5275 14170
rect 5327 14118 5339 14170
rect 5391 14118 12029 14170
rect 12081 14118 12093 14170
rect 12145 14118 12157 14170
rect 12209 14118 12221 14170
rect 12273 14118 12285 14170
rect 12337 14118 18975 14170
rect 19027 14118 19039 14170
rect 19091 14118 19103 14170
rect 19155 14118 19167 14170
rect 19219 14118 19231 14170
rect 19283 14118 25921 14170
rect 25973 14118 25985 14170
rect 26037 14118 26049 14170
rect 26101 14118 26113 14170
rect 26165 14118 26177 14170
rect 26229 14118 28888 14170
rect 1104 14096 28888 14118
rect 1104 13626 28888 13648
rect 1104 13574 4423 13626
rect 4475 13574 4487 13626
rect 4539 13574 4551 13626
rect 4603 13574 4615 13626
rect 4667 13574 4679 13626
rect 4731 13574 11369 13626
rect 11421 13574 11433 13626
rect 11485 13574 11497 13626
rect 11549 13574 11561 13626
rect 11613 13574 11625 13626
rect 11677 13574 18315 13626
rect 18367 13574 18379 13626
rect 18431 13574 18443 13626
rect 18495 13574 18507 13626
rect 18559 13574 18571 13626
rect 18623 13574 25261 13626
rect 25313 13574 25325 13626
rect 25377 13574 25389 13626
rect 25441 13574 25453 13626
rect 25505 13574 25517 13626
rect 25569 13574 28888 13626
rect 1104 13552 28888 13574
rect 16666 13268 16672 13320
rect 16724 13268 16730 13320
rect 16022 13132 16028 13184
rect 16080 13132 16086 13184
rect 1104 13082 28888 13104
rect 1104 13030 5083 13082
rect 5135 13030 5147 13082
rect 5199 13030 5211 13082
rect 5263 13030 5275 13082
rect 5327 13030 5339 13082
rect 5391 13030 12029 13082
rect 12081 13030 12093 13082
rect 12145 13030 12157 13082
rect 12209 13030 12221 13082
rect 12273 13030 12285 13082
rect 12337 13030 18975 13082
rect 19027 13030 19039 13082
rect 19091 13030 19103 13082
rect 19155 13030 19167 13082
rect 19219 13030 19231 13082
rect 19283 13030 25921 13082
rect 25973 13030 25985 13082
rect 26037 13030 26049 13082
rect 26101 13030 26113 13082
rect 26165 13030 26177 13082
rect 26229 13030 28888 13082
rect 1104 13008 28888 13030
rect 15838 12928 15844 12980
rect 15896 12928 15902 12980
rect 15933 12971 15991 12977
rect 15933 12937 15945 12971
rect 15979 12968 15991 12971
rect 16022 12968 16028 12980
rect 15979 12940 16028 12968
rect 15979 12937 15991 12940
rect 15933 12931 15991 12937
rect 16022 12928 16028 12940
rect 16080 12928 16086 12980
rect 15856 12900 15884 12928
rect 17037 12903 17095 12909
rect 15856 12872 16988 12900
rect 16485 12835 16543 12841
rect 16485 12801 16497 12835
rect 16531 12832 16543 12835
rect 16531 12804 16712 12832
rect 16531 12801 16543 12804
rect 16485 12795 16543 12801
rect 16117 12767 16175 12773
rect 16117 12733 16129 12767
rect 16163 12764 16175 12767
rect 16163 12736 16620 12764
rect 16163 12733 16175 12736
rect 16117 12727 16175 12733
rect 15470 12588 15476 12640
rect 15528 12588 15534 12640
rect 16298 12588 16304 12640
rect 16356 12588 16362 12640
rect 16592 12628 16620 12736
rect 16684 12705 16712 12804
rect 16669 12699 16727 12705
rect 16669 12665 16681 12699
rect 16715 12665 16727 12699
rect 16960 12696 16988 12872
rect 17037 12869 17049 12903
rect 17083 12900 17095 12903
rect 28258 12900 28264 12912
rect 17083 12872 28264 12900
rect 17083 12869 17095 12872
rect 17037 12863 17095 12869
rect 18432 12841 18460 12872
rect 28258 12860 28264 12872
rect 28316 12860 28322 12912
rect 17129 12835 17187 12841
rect 17129 12801 17141 12835
rect 17175 12832 17187 12835
rect 17497 12835 17555 12841
rect 17497 12832 17509 12835
rect 17175 12804 17509 12832
rect 17175 12801 17187 12804
rect 17129 12795 17187 12801
rect 17497 12801 17509 12804
rect 17543 12801 17555 12835
rect 17497 12795 17555 12801
rect 18417 12835 18475 12841
rect 18417 12801 18429 12835
rect 18463 12801 18475 12835
rect 18417 12795 18475 12801
rect 19242 12792 19248 12844
rect 19300 12792 19306 12844
rect 17310 12724 17316 12776
rect 17368 12724 17374 12776
rect 17402 12724 17408 12776
rect 17460 12764 17466 12776
rect 18049 12767 18107 12773
rect 18049 12764 18061 12767
rect 17460 12736 18061 12764
rect 17460 12724 17466 12736
rect 18049 12733 18061 12736
rect 18095 12733 18107 12767
rect 18049 12727 18107 12733
rect 18325 12767 18383 12773
rect 18325 12733 18337 12767
rect 18371 12733 18383 12767
rect 19153 12767 19211 12773
rect 19153 12764 19165 12767
rect 18325 12727 18383 12733
rect 18800 12736 19165 12764
rect 18340 12696 18368 12727
rect 18800 12705 18828 12736
rect 19153 12733 19165 12736
rect 19199 12733 19211 12767
rect 19153 12727 19211 12733
rect 16960 12668 18368 12696
rect 18785 12699 18843 12705
rect 16669 12659 16727 12665
rect 18785 12665 18797 12699
rect 18831 12665 18843 12699
rect 18785 12659 18843 12665
rect 18874 12656 18880 12708
rect 18932 12656 18938 12708
rect 17310 12628 17316 12640
rect 16592 12600 17316 12628
rect 17310 12588 17316 12600
rect 17368 12588 17374 12640
rect 1104 12538 28888 12560
rect 1104 12486 4423 12538
rect 4475 12486 4487 12538
rect 4539 12486 4551 12538
rect 4603 12486 4615 12538
rect 4667 12486 4679 12538
rect 4731 12486 11369 12538
rect 11421 12486 11433 12538
rect 11485 12486 11497 12538
rect 11549 12486 11561 12538
rect 11613 12486 11625 12538
rect 11677 12486 18315 12538
rect 18367 12486 18379 12538
rect 18431 12486 18443 12538
rect 18495 12486 18507 12538
rect 18559 12486 18571 12538
rect 18623 12486 25261 12538
rect 25313 12486 25325 12538
rect 25377 12486 25389 12538
rect 25441 12486 25453 12538
rect 25505 12486 25517 12538
rect 25569 12486 28888 12538
rect 1104 12464 28888 12486
rect 18141 12359 18199 12365
rect 18141 12325 18153 12359
rect 18187 12356 18199 12359
rect 19242 12356 19248 12368
rect 18187 12328 19248 12356
rect 18187 12325 18199 12328
rect 18141 12319 18199 12325
rect 19242 12316 19248 12328
rect 19300 12316 19306 12368
rect 15933 12291 15991 12297
rect 15933 12257 15945 12291
rect 15979 12288 15991 12291
rect 16298 12288 16304 12300
rect 15979 12260 16304 12288
rect 15979 12257 15991 12260
rect 15933 12251 15991 12257
rect 16298 12248 16304 12260
rect 16356 12248 16362 12300
rect 17865 12291 17923 12297
rect 17865 12257 17877 12291
rect 17911 12288 17923 12291
rect 17954 12288 17960 12300
rect 17911 12260 17960 12288
rect 17911 12257 17923 12260
rect 17865 12251 17923 12257
rect 17954 12248 17960 12260
rect 18012 12248 18018 12300
rect 15105 12223 15163 12229
rect 15105 12189 15117 12223
rect 15151 12220 15163 12223
rect 15470 12220 15476 12232
rect 15151 12192 15476 12220
rect 15151 12189 15163 12192
rect 15105 12183 15163 12189
rect 15470 12180 15476 12192
rect 15528 12180 15534 12232
rect 15657 12223 15715 12229
rect 15657 12189 15669 12223
rect 15703 12189 15715 12223
rect 15657 12183 15715 12189
rect 15672 12152 15700 12183
rect 17586 12180 17592 12232
rect 17644 12220 17650 12232
rect 17773 12223 17831 12229
rect 17773 12220 17785 12223
rect 17644 12192 17785 12220
rect 17644 12180 17650 12192
rect 17773 12189 17785 12192
rect 17819 12189 17831 12223
rect 17773 12183 17831 12189
rect 15120 12124 15700 12152
rect 15120 12096 15148 12124
rect 16482 12112 16488 12164
rect 16540 12112 16546 12164
rect 14918 12044 14924 12096
rect 14976 12044 14982 12096
rect 15102 12044 15108 12096
rect 15160 12044 15166 12096
rect 17402 12044 17408 12096
rect 17460 12044 17466 12096
rect 1104 11994 28888 12016
rect 1104 11942 5083 11994
rect 5135 11942 5147 11994
rect 5199 11942 5211 11994
rect 5263 11942 5275 11994
rect 5327 11942 5339 11994
rect 5391 11942 12029 11994
rect 12081 11942 12093 11994
rect 12145 11942 12157 11994
rect 12209 11942 12221 11994
rect 12273 11942 12285 11994
rect 12337 11942 18975 11994
rect 19027 11942 19039 11994
rect 19091 11942 19103 11994
rect 19155 11942 19167 11994
rect 19219 11942 19231 11994
rect 19283 11942 25921 11994
rect 25973 11942 25985 11994
rect 26037 11942 26049 11994
rect 26101 11942 26113 11994
rect 26165 11942 26177 11994
rect 26229 11942 28888 11994
rect 1104 11920 28888 11942
rect 14918 11840 14924 11892
rect 14976 11840 14982 11892
rect 17586 11840 17592 11892
rect 17644 11840 17650 11892
rect 14645 11815 14703 11821
rect 14645 11781 14657 11815
rect 14691 11812 14703 11815
rect 14936 11812 14964 11840
rect 21726 11812 21732 11824
rect 14691 11784 14964 11812
rect 21206 11784 21732 11812
rect 14691 11781 14703 11784
rect 14645 11775 14703 11781
rect 21726 11772 21732 11784
rect 21784 11772 21790 11824
rect 16482 11744 16488 11756
rect 15778 11716 16488 11744
rect 16482 11704 16488 11716
rect 16540 11704 16546 11756
rect 17681 11747 17739 11753
rect 17681 11713 17693 11747
rect 17727 11744 17739 11747
rect 18049 11747 18107 11753
rect 18049 11744 18061 11747
rect 17727 11716 18061 11744
rect 17727 11713 17739 11716
rect 17681 11707 17739 11713
rect 18049 11713 18061 11716
rect 18095 11713 18107 11747
rect 18049 11707 18107 11713
rect 18966 11704 18972 11756
rect 19024 11704 19030 11756
rect 19242 11704 19248 11756
rect 19300 11744 19306 11756
rect 19613 11747 19671 11753
rect 19613 11744 19625 11747
rect 19300 11716 19625 11744
rect 19300 11704 19306 11716
rect 19613 11713 19625 11716
rect 19659 11713 19671 11747
rect 19613 11707 19671 11713
rect 14369 11679 14427 11685
rect 14369 11645 14381 11679
rect 14415 11645 14427 11679
rect 14369 11639 14427 11645
rect 14182 11500 14188 11552
rect 14240 11540 14246 11552
rect 14384 11540 14412 11639
rect 17310 11636 17316 11688
rect 17368 11676 17374 11688
rect 17770 11676 17776 11688
rect 17368 11648 17776 11676
rect 17368 11636 17374 11648
rect 17770 11636 17776 11648
rect 17828 11636 17834 11688
rect 18601 11679 18659 11685
rect 18601 11676 18613 11679
rect 18064 11648 18613 11676
rect 16117 11611 16175 11617
rect 16117 11577 16129 11611
rect 16163 11608 16175 11611
rect 16666 11608 16672 11620
rect 16163 11580 16672 11608
rect 16163 11577 16175 11580
rect 16117 11571 16175 11577
rect 16666 11568 16672 11580
rect 16724 11608 16730 11620
rect 16724 11580 17540 11608
rect 16724 11568 16730 11580
rect 17512 11552 17540 11580
rect 18064 11552 18092 11648
rect 18601 11645 18613 11648
rect 18647 11645 18659 11679
rect 18601 11639 18659 11645
rect 18877 11679 18935 11685
rect 18877 11645 18889 11679
rect 18923 11645 18935 11679
rect 18877 11639 18935 11645
rect 19797 11679 19855 11685
rect 19797 11645 19809 11679
rect 19843 11676 19855 11679
rect 19978 11676 19984 11688
rect 19843 11648 19984 11676
rect 19843 11645 19855 11648
rect 19797 11639 19855 11645
rect 18230 11568 18236 11620
rect 18288 11608 18294 11620
rect 18892 11608 18920 11639
rect 19978 11636 19984 11648
rect 20036 11636 20042 11688
rect 20162 11636 20168 11688
rect 20220 11636 20226 11688
rect 18288 11580 18920 11608
rect 18288 11568 18294 11580
rect 19334 11568 19340 11620
rect 19392 11568 19398 11620
rect 15102 11540 15108 11552
rect 14240 11512 15108 11540
rect 14240 11500 14246 11512
rect 15102 11500 15108 11512
rect 15160 11500 15166 11552
rect 17218 11500 17224 11552
rect 17276 11500 17282 11552
rect 17494 11500 17500 11552
rect 17552 11500 17558 11552
rect 18046 11500 18052 11552
rect 18104 11500 18110 11552
rect 19426 11500 19432 11552
rect 19484 11500 19490 11552
rect 21634 11549 21640 11552
rect 21591 11543 21640 11549
rect 21591 11509 21603 11543
rect 21637 11509 21640 11543
rect 21591 11503 21640 11509
rect 21634 11500 21640 11503
rect 21692 11500 21698 11552
rect 1104 11450 28888 11472
rect 1104 11398 4423 11450
rect 4475 11398 4487 11450
rect 4539 11398 4551 11450
rect 4603 11398 4615 11450
rect 4667 11398 4679 11450
rect 4731 11398 11369 11450
rect 11421 11398 11433 11450
rect 11485 11398 11497 11450
rect 11549 11398 11561 11450
rect 11613 11398 11625 11450
rect 11677 11398 18315 11450
rect 18367 11398 18379 11450
rect 18431 11398 18443 11450
rect 18495 11398 18507 11450
rect 18559 11398 18571 11450
rect 18623 11398 25261 11450
rect 25313 11398 25325 11450
rect 25377 11398 25389 11450
rect 25441 11398 25453 11450
rect 25505 11398 25517 11450
rect 25569 11398 28888 11450
rect 1104 11376 28888 11398
rect 13817 11339 13875 11345
rect 13817 11305 13829 11339
rect 13863 11336 13875 11339
rect 16574 11336 16580 11348
rect 13863 11308 16580 11336
rect 13863 11305 13875 11308
rect 13817 11299 13875 11305
rect 16574 11296 16580 11308
rect 16632 11296 16638 11348
rect 19242 11296 19248 11348
rect 19300 11296 19306 11348
rect 20990 11296 20996 11348
rect 21048 11336 21054 11348
rect 21450 11336 21456 11348
rect 21048 11308 21456 11336
rect 21048 11296 21054 11308
rect 21450 11296 21456 11308
rect 21508 11296 21514 11348
rect 17957 11271 18015 11277
rect 17957 11237 17969 11271
rect 18003 11268 18015 11271
rect 18046 11268 18052 11280
rect 18003 11240 18052 11268
rect 18003 11237 18015 11240
rect 17957 11231 18015 11237
rect 18046 11228 18052 11240
rect 18104 11228 18110 11280
rect 13446 11160 13452 11212
rect 13504 11200 13510 11212
rect 13814 11200 13820 11212
rect 13504 11172 13820 11200
rect 13504 11160 13510 11172
rect 13814 11160 13820 11172
rect 13872 11160 13878 11212
rect 14461 11203 14519 11209
rect 14461 11169 14473 11203
rect 14507 11200 14519 11203
rect 15010 11200 15016 11212
rect 14507 11172 15016 11200
rect 14507 11169 14519 11172
rect 14461 11163 14519 11169
rect 15010 11160 15016 11172
rect 15068 11160 15074 11212
rect 16482 11200 16488 11212
rect 15764 11172 16488 11200
rect 13538 11092 13544 11144
rect 13596 11092 13602 11144
rect 14182 11092 14188 11144
rect 14240 11092 14246 11144
rect 15764 11076 15792 11172
rect 16482 11160 16488 11172
rect 16540 11200 16546 11212
rect 16540 11172 17724 11200
rect 16540 11160 16546 11172
rect 16209 11135 16267 11141
rect 16209 11101 16221 11135
rect 16255 11101 16267 11135
rect 16209 11095 16267 11101
rect 15746 11064 15752 11076
rect 15686 11036 15752 11064
rect 15746 11024 15752 11036
rect 15804 11024 15810 11076
rect 16224 11064 16252 11095
rect 16485 11067 16543 11073
rect 16224 11036 16344 11064
rect 16316 11008 16344 11036
rect 16485 11033 16497 11067
rect 16531 11064 16543 11067
rect 17696 11064 17724 11172
rect 17770 11160 17776 11212
rect 17828 11200 17834 11212
rect 19797 11203 19855 11209
rect 19797 11200 19809 11203
rect 17828 11172 19809 11200
rect 17828 11160 17834 11172
rect 19797 11169 19809 11172
rect 19843 11169 19855 11203
rect 19797 11163 19855 11169
rect 18782 11092 18788 11144
rect 18840 11132 18846 11144
rect 18969 11135 19027 11141
rect 18969 11132 18981 11135
rect 18840 11104 18981 11132
rect 18840 11092 18846 11104
rect 18969 11101 18981 11104
rect 19015 11101 19027 11135
rect 18969 11095 19027 11101
rect 19334 11092 19340 11144
rect 19392 11132 19398 11144
rect 19613 11135 19671 11141
rect 19613 11132 19625 11135
rect 19392 11104 19625 11132
rect 19392 11092 19398 11104
rect 19613 11101 19625 11104
rect 19659 11101 19671 11135
rect 19613 11095 19671 11101
rect 20714 11092 20720 11144
rect 20772 11092 20778 11144
rect 22741 11135 22799 11141
rect 22741 11101 22753 11135
rect 22787 11101 22799 11135
rect 22741 11095 22799 11101
rect 19705 11067 19763 11073
rect 16531 11036 16896 11064
rect 17696 11050 18552 11064
rect 17710 11036 18552 11050
rect 16531 11033 16543 11036
rect 16485 11027 16543 11033
rect 15930 10956 15936 11008
rect 15988 10956 15994 11008
rect 16298 10956 16304 11008
rect 16356 10956 16362 11008
rect 16868 10996 16896 11036
rect 17310 10996 17316 11008
rect 16868 10968 17316 10996
rect 17310 10956 17316 10968
rect 17368 10956 17374 11008
rect 18138 10956 18144 11008
rect 18196 10996 18202 11008
rect 18417 10999 18475 11005
rect 18417 10996 18429 10999
rect 18196 10968 18429 10996
rect 18196 10956 18202 10968
rect 18417 10965 18429 10968
rect 18463 10965 18475 10999
rect 18524 10996 18552 11036
rect 19705 11033 19717 11067
rect 19751 11064 19763 11067
rect 20073 11067 20131 11073
rect 20073 11064 20085 11067
rect 19751 11036 20085 11064
rect 19751 11033 19763 11036
rect 19705 11027 19763 11033
rect 20073 11033 20085 11036
rect 20119 11033 20131 11067
rect 20073 11027 20131 11033
rect 22002 11024 22008 11076
rect 22060 11024 22066 11076
rect 22462 11024 22468 11076
rect 22520 11024 22526 11076
rect 22756 11064 22784 11095
rect 22572 11036 22784 11064
rect 22572 11008 22600 11036
rect 18874 10996 18880 11008
rect 18524 10968 18880 10996
rect 18417 10959 18475 10965
rect 18874 10956 18880 10968
rect 18932 10956 18938 11008
rect 22554 10956 22560 11008
rect 22612 10956 22618 11008
rect 1104 10906 28888 10928
rect 1104 10854 5083 10906
rect 5135 10854 5147 10906
rect 5199 10854 5211 10906
rect 5263 10854 5275 10906
rect 5327 10854 5339 10906
rect 5391 10854 12029 10906
rect 12081 10854 12093 10906
rect 12145 10854 12157 10906
rect 12209 10854 12221 10906
rect 12273 10854 12285 10906
rect 12337 10854 18975 10906
rect 19027 10854 19039 10906
rect 19091 10854 19103 10906
rect 19155 10854 19167 10906
rect 19219 10854 19231 10906
rect 19283 10854 25921 10906
rect 25973 10854 25985 10906
rect 26037 10854 26049 10906
rect 26101 10854 26113 10906
rect 26165 10854 26177 10906
rect 26229 10854 28888 10906
rect 1104 10832 28888 10854
rect 13814 10752 13820 10804
rect 13872 10792 13878 10804
rect 14553 10795 14611 10801
rect 14553 10792 14565 10795
rect 13872 10764 14565 10792
rect 13872 10752 13878 10764
rect 14553 10761 14565 10764
rect 14599 10761 14611 10795
rect 14553 10755 14611 10761
rect 14921 10795 14979 10801
rect 14921 10761 14933 10795
rect 14967 10761 14979 10795
rect 14921 10755 14979 10761
rect 14936 10656 14964 10755
rect 15010 10752 15016 10804
rect 15068 10752 15074 10804
rect 17218 10752 17224 10804
rect 17276 10752 17282 10804
rect 17310 10752 17316 10804
rect 17368 10752 17374 10804
rect 17865 10795 17923 10801
rect 17865 10761 17877 10795
rect 17911 10792 17923 10795
rect 18138 10792 18144 10804
rect 17911 10764 18144 10792
rect 17911 10761 17923 10764
rect 17865 10755 17923 10761
rect 18138 10752 18144 10764
rect 18196 10752 18202 10804
rect 18325 10795 18383 10801
rect 18325 10761 18337 10795
rect 18371 10761 18383 10795
rect 18325 10755 18383 10761
rect 20441 10795 20499 10801
rect 20441 10761 20453 10795
rect 20487 10792 20499 10795
rect 20714 10792 20720 10804
rect 20487 10764 20720 10792
rect 20487 10761 20499 10764
rect 20441 10755 20499 10761
rect 15197 10659 15255 10665
rect 15197 10656 15209 10659
rect 14936 10628 15209 10656
rect 15197 10625 15209 10628
rect 15243 10625 15255 10659
rect 15197 10619 15255 10625
rect 16390 10616 16396 10668
rect 16448 10656 16454 10668
rect 16853 10659 16911 10665
rect 16853 10656 16865 10659
rect 16448 10628 16865 10656
rect 16448 10616 16454 10628
rect 16853 10625 16865 10628
rect 16899 10625 16911 10659
rect 17236 10656 17264 10752
rect 17497 10659 17555 10665
rect 17497 10656 17509 10659
rect 17236 10628 17509 10656
rect 16853 10619 16911 10625
rect 17497 10625 17509 10628
rect 17543 10625 17555 10659
rect 17497 10619 17555 10625
rect 17954 10616 17960 10668
rect 18012 10616 18018 10668
rect 18340 10656 18368 10755
rect 20714 10752 20720 10764
rect 20772 10752 20778 10804
rect 21453 10795 21511 10801
rect 21453 10761 21465 10795
rect 21499 10792 21511 10795
rect 22462 10792 22468 10804
rect 21499 10764 22468 10792
rect 21499 10761 21511 10764
rect 21453 10755 21511 10761
rect 22462 10752 22468 10764
rect 22520 10752 22526 10804
rect 23934 10792 23940 10804
rect 23308 10764 23940 10792
rect 19702 10684 19708 10736
rect 19760 10684 19766 10736
rect 23308 10724 23336 10764
rect 23934 10752 23940 10764
rect 23992 10792 23998 10804
rect 23992 10764 24716 10792
rect 23992 10752 23998 10764
rect 24688 10733 24716 10764
rect 22066 10696 23336 10724
rect 24673 10727 24731 10733
rect 18601 10659 18659 10665
rect 18601 10656 18613 10659
rect 18340 10628 18613 10656
rect 18601 10625 18613 10628
rect 18647 10625 18659 10659
rect 18601 10619 18659 10625
rect 21266 10616 21272 10668
rect 21324 10616 21330 10668
rect 21818 10616 21824 10668
rect 21876 10656 21882 10668
rect 21913 10659 21971 10665
rect 21913 10656 21925 10659
rect 21876 10628 21925 10656
rect 21876 10616 21882 10628
rect 21913 10625 21925 10628
rect 21959 10656 21971 10659
rect 22066 10656 22094 10696
rect 24673 10693 24685 10727
rect 24719 10693 24731 10727
rect 24673 10687 24731 10693
rect 21959 10628 22094 10656
rect 22189 10659 22247 10665
rect 21959 10625 21971 10628
rect 21913 10619 21971 10625
rect 22189 10625 22201 10659
rect 22235 10625 22247 10659
rect 22189 10619 22247 10625
rect 14369 10591 14427 10597
rect 14369 10557 14381 10591
rect 14415 10557 14427 10591
rect 14369 10551 14427 10557
rect 14461 10591 14519 10597
rect 14461 10557 14473 10591
rect 14507 10588 14519 10591
rect 15289 10591 15347 10597
rect 15289 10588 15301 10591
rect 14507 10560 15301 10588
rect 14507 10557 14519 10560
rect 14461 10551 14519 10557
rect 15289 10557 15301 10560
rect 15335 10557 15347 10591
rect 15289 10551 15347 10557
rect 14384 10520 14412 10551
rect 15930 10548 15936 10600
rect 15988 10588 15994 10600
rect 16482 10588 16488 10600
rect 15988 10560 16488 10588
rect 15988 10548 15994 10560
rect 16482 10548 16488 10560
rect 16540 10548 16546 10600
rect 16574 10548 16580 10600
rect 16632 10588 16638 10600
rect 16761 10591 16819 10597
rect 16761 10588 16773 10591
rect 16632 10560 16773 10588
rect 16632 10548 16638 10560
rect 16761 10557 16773 10560
rect 16807 10557 16819 10591
rect 16761 10551 16819 10557
rect 17770 10548 17776 10600
rect 17828 10548 17834 10600
rect 18230 10548 18236 10600
rect 18288 10548 18294 10600
rect 18693 10591 18751 10597
rect 18693 10557 18705 10591
rect 18739 10557 18751 10591
rect 18693 10551 18751 10557
rect 18969 10591 19027 10597
rect 18969 10557 18981 10591
rect 19015 10588 19027 10591
rect 19426 10588 19432 10600
rect 19015 10560 19432 10588
rect 19015 10557 19027 10560
rect 18969 10551 19027 10557
rect 17221 10523 17279 10529
rect 14384 10492 15056 10520
rect 15028 10464 15056 10492
rect 17221 10489 17233 10523
rect 17267 10520 17279 10523
rect 18248 10520 18276 10548
rect 17267 10492 18276 10520
rect 17267 10489 17279 10492
rect 17221 10483 17279 10489
rect 18708 10464 18736 10551
rect 19426 10548 19432 10560
rect 19484 10548 19490 10600
rect 21910 10480 21916 10532
rect 21968 10480 21974 10532
rect 15010 10412 15016 10464
rect 15068 10412 15074 10464
rect 18230 10412 18236 10464
rect 18288 10452 18294 10464
rect 18417 10455 18475 10461
rect 18417 10452 18429 10455
rect 18288 10424 18429 10452
rect 18288 10412 18294 10424
rect 18417 10421 18429 10424
rect 18463 10421 18475 10455
rect 18417 10415 18475 10421
rect 18690 10412 18696 10464
rect 18748 10452 18754 10464
rect 19978 10452 19984 10464
rect 18748 10424 19984 10452
rect 18748 10412 18754 10424
rect 19978 10412 19984 10424
rect 20036 10412 20042 10464
rect 21542 10412 21548 10464
rect 21600 10452 21606 10464
rect 22204 10452 22232 10619
rect 22278 10616 22284 10668
rect 22336 10616 22342 10668
rect 24026 10616 24032 10668
rect 24084 10616 24090 10668
rect 22554 10548 22560 10600
rect 22612 10588 22618 10600
rect 22649 10591 22707 10597
rect 22649 10588 22661 10591
rect 22612 10560 22661 10588
rect 22612 10548 22618 10560
rect 22649 10557 22661 10560
rect 22695 10557 22707 10591
rect 22925 10591 22983 10597
rect 22925 10588 22937 10591
rect 22649 10551 22707 10557
rect 22756 10560 22937 10588
rect 22465 10523 22523 10529
rect 22465 10489 22477 10523
rect 22511 10520 22523 10523
rect 22756 10520 22784 10560
rect 22925 10557 22937 10560
rect 22971 10557 22983 10591
rect 22925 10551 22983 10557
rect 22511 10492 22784 10520
rect 22511 10489 22523 10492
rect 22465 10483 22523 10489
rect 24302 10452 24308 10464
rect 21600 10424 24308 10452
rect 21600 10412 21606 10424
rect 24302 10412 24308 10424
rect 24360 10412 24366 10464
rect 1104 10362 28888 10384
rect 1104 10310 4423 10362
rect 4475 10310 4487 10362
rect 4539 10310 4551 10362
rect 4603 10310 4615 10362
rect 4667 10310 4679 10362
rect 4731 10310 11369 10362
rect 11421 10310 11433 10362
rect 11485 10310 11497 10362
rect 11549 10310 11561 10362
rect 11613 10310 11625 10362
rect 11677 10310 18315 10362
rect 18367 10310 18379 10362
rect 18431 10310 18443 10362
rect 18495 10310 18507 10362
rect 18559 10310 18571 10362
rect 18623 10310 25261 10362
rect 25313 10310 25325 10362
rect 25377 10310 25389 10362
rect 25441 10310 25453 10362
rect 25505 10310 25517 10362
rect 25569 10310 28888 10362
rect 1104 10288 28888 10310
rect 15102 10248 15108 10260
rect 14108 10220 15108 10248
rect 14108 10121 14136 10220
rect 15102 10208 15108 10220
rect 15160 10248 15166 10260
rect 16298 10248 16304 10260
rect 15160 10220 16304 10248
rect 15160 10208 15166 10220
rect 16298 10208 16304 10220
rect 16356 10248 16362 10260
rect 18690 10248 18696 10260
rect 16356 10220 18696 10248
rect 16356 10208 16362 10220
rect 16960 10121 16988 10220
rect 18690 10208 18696 10220
rect 18748 10208 18754 10260
rect 18782 10208 18788 10260
rect 18840 10208 18846 10260
rect 20806 10208 20812 10260
rect 20864 10248 20870 10260
rect 22002 10248 22008 10260
rect 20864 10220 22008 10248
rect 20864 10208 20870 10220
rect 22002 10208 22008 10220
rect 22060 10248 22066 10260
rect 22060 10220 23704 10248
rect 22060 10208 22066 10220
rect 18230 10140 18236 10192
rect 18288 10140 18294 10192
rect 14093 10115 14151 10121
rect 14093 10081 14105 10115
rect 14139 10081 14151 10115
rect 14093 10075 14151 10081
rect 16945 10115 17003 10121
rect 16945 10081 16957 10115
rect 16991 10081 17003 10115
rect 16945 10075 17003 10081
rect 17221 10115 17279 10121
rect 17221 10081 17233 10115
rect 17267 10112 17279 10115
rect 18248 10112 18276 10140
rect 17267 10084 18276 10112
rect 18693 10115 18751 10121
rect 17267 10081 17279 10084
rect 17221 10075 17279 10081
rect 18693 10081 18705 10115
rect 18739 10112 18751 10115
rect 18800 10112 18828 10208
rect 21358 10180 21364 10192
rect 18739 10084 18828 10112
rect 20088 10152 21364 10180
rect 18739 10081 18751 10084
rect 18693 10075 18751 10081
rect 15746 10044 15752 10056
rect 15502 10016 15752 10044
rect 15746 10004 15752 10016
rect 15804 10004 15810 10056
rect 20088 10053 20116 10152
rect 21358 10140 21364 10152
rect 21416 10140 21422 10192
rect 20533 10115 20591 10121
rect 20533 10081 20545 10115
rect 20579 10112 20591 10115
rect 20714 10112 20720 10124
rect 20579 10084 20720 10112
rect 20579 10081 20591 10084
rect 20533 10075 20591 10081
rect 20714 10072 20720 10084
rect 20772 10072 20778 10124
rect 21545 10115 21603 10121
rect 21100 10084 21496 10112
rect 21100 10056 21128 10084
rect 16577 10047 16635 10053
rect 16577 10013 16589 10047
rect 16623 10013 16635 10047
rect 16577 10007 16635 10013
rect 20073 10047 20131 10053
rect 20073 10013 20085 10047
rect 20119 10013 20131 10047
rect 20073 10007 20131 10013
rect 14366 9936 14372 9988
rect 14424 9936 14430 9988
rect 16592 9976 16620 10007
rect 21082 10004 21088 10056
rect 21140 10004 21146 10056
rect 21174 10004 21180 10056
rect 21232 10004 21238 10056
rect 21468 10044 21496 10084
rect 21545 10081 21557 10115
rect 21591 10112 21603 10115
rect 21634 10112 21640 10124
rect 21591 10084 21640 10112
rect 21591 10081 21603 10084
rect 21545 10075 21603 10081
rect 21634 10072 21640 10084
rect 21692 10072 21698 10124
rect 22189 10115 22247 10121
rect 22189 10081 22201 10115
rect 22235 10112 22247 10115
rect 22554 10112 22560 10124
rect 22235 10084 22560 10112
rect 22235 10081 22247 10084
rect 22189 10075 22247 10081
rect 22554 10072 22560 10084
rect 22612 10112 22618 10124
rect 23198 10112 23204 10124
rect 22612 10084 23204 10112
rect 22612 10072 22618 10084
rect 23198 10072 23204 10084
rect 23256 10072 23262 10124
rect 21818 10044 21824 10056
rect 21468 10016 21824 10044
rect 21818 10004 21824 10016
rect 21876 10004 21882 10056
rect 22002 10004 22008 10056
rect 22060 10004 22066 10056
rect 18690 9976 18696 9988
rect 15856 9948 17632 9976
rect 18446 9948 18696 9976
rect 15856 9917 15884 9948
rect 17604 9920 17632 9948
rect 18690 9936 18696 9948
rect 18748 9976 18754 9988
rect 18874 9976 18880 9988
rect 18748 9948 18880 9976
rect 18748 9936 18754 9948
rect 18874 9936 18880 9948
rect 18932 9936 18938 9988
rect 19610 9936 19616 9988
rect 19668 9976 19674 9988
rect 20165 9979 20223 9985
rect 20165 9976 20177 9979
rect 19668 9948 20177 9976
rect 19668 9936 19674 9948
rect 20165 9945 20177 9948
rect 20211 9945 20223 9979
rect 20165 9939 20223 9945
rect 20254 9936 20260 9988
rect 20312 9936 20318 9988
rect 20395 9979 20453 9985
rect 20395 9945 20407 9979
rect 20441 9976 20453 9979
rect 21453 9979 21511 9985
rect 20441 9948 21404 9976
rect 20441 9945 20453 9948
rect 20395 9939 20453 9945
rect 15841 9911 15899 9917
rect 15841 9877 15853 9911
rect 15887 9877 15899 9911
rect 15841 9871 15899 9877
rect 15930 9868 15936 9920
rect 15988 9868 15994 9920
rect 17586 9868 17592 9920
rect 17644 9868 17650 9920
rect 19889 9911 19947 9917
rect 19889 9877 19901 9911
rect 19935 9908 19947 9911
rect 20530 9908 20536 9920
rect 19935 9880 20536 9908
rect 19935 9877 19947 9880
rect 19889 9871 19947 9877
rect 20530 9868 20536 9880
rect 20588 9868 20594 9920
rect 20898 9868 20904 9920
rect 20956 9868 20962 9920
rect 21376 9908 21404 9948
rect 21453 9945 21465 9979
rect 21499 9976 21511 9979
rect 21542 9976 21548 9988
rect 21499 9948 21548 9976
rect 21499 9945 21511 9948
rect 21453 9939 21511 9945
rect 21542 9936 21548 9948
rect 21600 9936 21606 9988
rect 22462 9936 22468 9988
rect 22520 9936 22526 9988
rect 23676 9976 23704 10220
rect 24026 9976 24032 9988
rect 23676 9962 24032 9976
rect 23690 9948 24032 9962
rect 24026 9936 24032 9948
rect 24084 9936 24090 9988
rect 24213 9979 24271 9985
rect 24213 9945 24225 9979
rect 24259 9976 24271 9979
rect 24302 9976 24308 9988
rect 24259 9948 24308 9976
rect 24259 9945 24271 9948
rect 24213 9939 24271 9945
rect 24302 9936 24308 9948
rect 24360 9936 24366 9988
rect 21637 9911 21695 9917
rect 21637 9908 21649 9911
rect 21376 9880 21649 9908
rect 21637 9877 21649 9880
rect 21683 9908 21695 9911
rect 22554 9908 22560 9920
rect 21683 9880 22560 9908
rect 21683 9877 21695 9880
rect 21637 9871 21695 9877
rect 22554 9868 22560 9880
rect 22612 9868 22618 9920
rect 1104 9818 28888 9840
rect 1104 9766 5083 9818
rect 5135 9766 5147 9818
rect 5199 9766 5211 9818
rect 5263 9766 5275 9818
rect 5327 9766 5339 9818
rect 5391 9766 12029 9818
rect 12081 9766 12093 9818
rect 12145 9766 12157 9818
rect 12209 9766 12221 9818
rect 12273 9766 12285 9818
rect 12337 9766 18975 9818
rect 19027 9766 19039 9818
rect 19091 9766 19103 9818
rect 19155 9766 19167 9818
rect 19219 9766 19231 9818
rect 19283 9766 25921 9818
rect 25973 9766 25985 9818
rect 26037 9766 26049 9818
rect 26101 9766 26113 9818
rect 26165 9766 26177 9818
rect 26229 9766 28888 9818
rect 1104 9744 28888 9766
rect 14366 9664 14372 9716
rect 14424 9704 14430 9716
rect 14921 9707 14979 9713
rect 14921 9704 14933 9707
rect 14424 9676 14933 9704
rect 14424 9664 14430 9676
rect 14921 9673 14933 9676
rect 14967 9673 14979 9707
rect 14921 9667 14979 9673
rect 15930 9664 15936 9716
rect 15988 9664 15994 9716
rect 19610 9664 19616 9716
rect 19668 9664 19674 9716
rect 20806 9704 20812 9716
rect 19720 9676 20812 9704
rect 15948 9636 15976 9664
rect 19720 9636 19748 9676
rect 20806 9664 20812 9676
rect 20864 9664 20870 9716
rect 21910 9664 21916 9716
rect 21968 9664 21974 9716
rect 22189 9707 22247 9713
rect 22189 9673 22201 9707
rect 22235 9704 22247 9707
rect 22278 9704 22284 9716
rect 22235 9676 22284 9704
rect 22235 9673 22247 9676
rect 22189 9667 22247 9673
rect 22278 9664 22284 9676
rect 22336 9664 22342 9716
rect 22462 9664 22468 9716
rect 22520 9704 22526 9716
rect 23017 9707 23075 9713
rect 23017 9704 23029 9707
rect 22520 9676 23029 9704
rect 22520 9664 22526 9676
rect 23017 9673 23029 9676
rect 23063 9673 23075 9707
rect 23017 9667 23075 9673
rect 21085 9639 21143 9645
rect 21085 9636 21097 9639
rect 14384 9608 15976 9636
rect 18892 9608 19748 9636
rect 19812 9608 21097 9636
rect 13538 9528 13544 9580
rect 13596 9568 13602 9580
rect 14384 9577 14412 9608
rect 14369 9571 14427 9577
rect 13596 9540 14320 9568
rect 13596 9528 13602 9540
rect 14185 9503 14243 9509
rect 14185 9469 14197 9503
rect 14231 9469 14243 9503
rect 14292 9500 14320 9540
rect 14369 9537 14381 9571
rect 14415 9537 14427 9571
rect 14369 9531 14427 9537
rect 14461 9571 14519 9577
rect 14461 9537 14473 9571
rect 14507 9537 14519 9571
rect 15105 9571 15163 9577
rect 15105 9568 15117 9571
rect 14461 9531 14519 9537
rect 14844 9540 15117 9568
rect 14476 9500 14504 9531
rect 14292 9472 14504 9500
rect 14185 9463 14243 9469
rect 14200 9432 14228 9463
rect 14734 9460 14740 9512
rect 14792 9460 14798 9512
rect 14752 9432 14780 9460
rect 14844 9441 14872 9540
rect 15105 9537 15117 9540
rect 15151 9537 15163 9571
rect 15105 9531 15163 9537
rect 15473 9571 15531 9577
rect 15473 9537 15485 9571
rect 15519 9537 15531 9571
rect 15473 9531 15531 9537
rect 14200 9404 14780 9432
rect 14829 9435 14887 9441
rect 14829 9401 14841 9435
rect 14875 9401 14887 9435
rect 14829 9395 14887 9401
rect 14734 9324 14740 9376
rect 14792 9364 14798 9376
rect 15488 9364 15516 9531
rect 17402 9528 17408 9580
rect 17460 9528 17466 9580
rect 18230 9528 18236 9580
rect 18288 9528 18294 9580
rect 18417 9571 18475 9577
rect 18417 9537 18429 9571
rect 18463 9568 18475 9571
rect 18782 9568 18788 9580
rect 18463 9540 18788 9568
rect 18463 9537 18475 9540
rect 18417 9531 18475 9537
rect 18782 9528 18788 9540
rect 18840 9528 18846 9580
rect 15565 9503 15623 9509
rect 15565 9469 15577 9503
rect 15611 9469 15623 9503
rect 15565 9463 15623 9469
rect 15841 9503 15899 9509
rect 15841 9469 15853 9503
rect 15887 9500 15899 9503
rect 16390 9500 16396 9512
rect 15887 9472 16396 9500
rect 15887 9469 15899 9472
rect 15841 9463 15899 9469
rect 15580 9432 15608 9463
rect 16390 9460 16396 9472
rect 16448 9460 16454 9512
rect 16482 9460 16488 9512
rect 16540 9500 16546 9512
rect 17543 9503 17601 9509
rect 17543 9500 17555 9503
rect 16540 9472 17555 9500
rect 16540 9460 16546 9472
rect 17543 9469 17555 9472
rect 17589 9469 17601 9503
rect 17543 9463 17601 9469
rect 17678 9460 17684 9512
rect 17736 9460 17742 9512
rect 18248 9500 18276 9528
rect 18601 9503 18659 9509
rect 18601 9500 18613 9503
rect 18248 9472 18613 9500
rect 18601 9469 18613 9472
rect 18647 9469 18659 9503
rect 18601 9463 18659 9469
rect 17957 9435 18015 9441
rect 15580 9404 16896 9432
rect 14792 9336 15516 9364
rect 14792 9324 14798 9336
rect 16758 9324 16764 9376
rect 16816 9324 16822 9376
rect 16868 9364 16896 9404
rect 17957 9401 17969 9435
rect 18003 9401 18015 9435
rect 17957 9395 18015 9401
rect 17218 9364 17224 9376
rect 16868 9336 17224 9364
rect 17218 9324 17224 9336
rect 17276 9324 17282 9376
rect 17310 9324 17316 9376
rect 17368 9364 17374 9376
rect 17678 9364 17684 9376
rect 17368 9336 17684 9364
rect 17368 9324 17374 9336
rect 17678 9324 17684 9336
rect 17736 9324 17742 9376
rect 17972 9364 18000 9395
rect 18138 9392 18144 9444
rect 18196 9432 18202 9444
rect 18782 9432 18788 9444
rect 18196 9404 18788 9432
rect 18196 9392 18202 9404
rect 18782 9392 18788 9404
rect 18840 9432 18846 9444
rect 18892 9432 18920 9608
rect 19812 9577 19840 9608
rect 21085 9605 21097 9608
rect 21131 9605 21143 9639
rect 21358 9636 21364 9648
rect 21085 9599 21143 9605
rect 21192 9608 21364 9636
rect 19153 9571 19211 9577
rect 19153 9537 19165 9571
rect 19199 9568 19211 9571
rect 19797 9571 19855 9577
rect 19199 9540 19380 9568
rect 19199 9537 19211 9540
rect 19153 9531 19211 9537
rect 18840 9404 18920 9432
rect 19352 9500 19380 9540
rect 19797 9537 19809 9571
rect 19843 9537 19855 9571
rect 19797 9531 19855 9537
rect 20809 9571 20867 9577
rect 20809 9537 20821 9571
rect 20855 9568 20867 9571
rect 20898 9568 20904 9580
rect 20855 9540 20904 9568
rect 20855 9537 20867 9540
rect 20809 9531 20867 9537
rect 20898 9528 20904 9540
rect 20956 9528 20962 9580
rect 20990 9528 20996 9580
rect 21048 9528 21054 9580
rect 21192 9577 21220 9608
rect 21358 9596 21364 9608
rect 21416 9636 21422 9648
rect 21928 9636 21956 9664
rect 21416 9608 21956 9636
rect 21416 9596 21422 9608
rect 22002 9596 22008 9648
rect 22060 9636 22066 9648
rect 22060 9608 23244 9636
rect 22060 9596 22066 9608
rect 21177 9571 21235 9577
rect 21177 9537 21189 9571
rect 21223 9537 21235 9571
rect 21177 9531 21235 9537
rect 21634 9528 21640 9580
rect 21692 9568 21698 9580
rect 21913 9571 21971 9577
rect 21913 9568 21925 9571
rect 21692 9540 21925 9568
rect 21692 9528 21698 9540
rect 21913 9537 21925 9540
rect 21959 9537 21971 9571
rect 21913 9531 21971 9537
rect 19889 9503 19947 9509
rect 19889 9500 19901 9503
rect 19352 9472 19901 9500
rect 18840 9392 18846 9404
rect 19352 9376 19380 9472
rect 19889 9469 19901 9472
rect 19935 9469 19947 9503
rect 19889 9463 19947 9469
rect 19981 9503 20039 9509
rect 19981 9469 19993 9503
rect 20027 9469 20039 9503
rect 19981 9463 20039 9469
rect 19426 9392 19432 9444
rect 19484 9432 19490 9444
rect 19996 9432 20024 9463
rect 20070 9460 20076 9512
rect 20128 9460 20134 9512
rect 20530 9460 20536 9512
rect 20588 9460 20594 9512
rect 22020 9509 22048 9596
rect 23216 9577 23244 9608
rect 22557 9571 22615 9577
rect 22557 9537 22569 9571
rect 22603 9537 22615 9571
rect 22557 9531 22615 9537
rect 23201 9571 23259 9577
rect 23201 9537 23213 9571
rect 23247 9537 23259 9571
rect 23201 9531 23259 9537
rect 23293 9571 23351 9577
rect 23293 9537 23305 9571
rect 23339 9537 23351 9571
rect 23293 9531 23351 9537
rect 23569 9571 23627 9577
rect 23569 9537 23581 9571
rect 23615 9568 23627 9571
rect 23615 9540 24164 9568
rect 23615 9537 23627 9540
rect 23569 9531 23627 9537
rect 20625 9503 20683 9509
rect 20625 9469 20637 9503
rect 20671 9469 20683 9503
rect 20625 9463 20683 9469
rect 20717 9503 20775 9509
rect 20717 9469 20729 9503
rect 20763 9500 20775 9503
rect 22005 9503 22063 9509
rect 22005 9500 22017 9503
rect 20763 9472 22017 9500
rect 20763 9469 20775 9472
rect 20717 9463 20775 9469
rect 22005 9469 22017 9472
rect 22051 9469 22063 9503
rect 22005 9463 22063 9469
rect 19484 9404 20024 9432
rect 19484 9392 19490 9404
rect 20162 9392 20168 9444
rect 20220 9432 20226 9444
rect 20349 9435 20407 9441
rect 20349 9432 20361 9435
rect 20220 9404 20361 9432
rect 20220 9392 20226 9404
rect 20349 9401 20361 9404
rect 20395 9401 20407 9435
rect 20640 9432 20668 9463
rect 20640 9404 21036 9432
rect 20349 9395 20407 9401
rect 21008 9376 21036 9404
rect 21082 9392 21088 9444
rect 21140 9432 21146 9444
rect 22572 9432 22600 9531
rect 22646 9460 22652 9512
rect 22704 9460 22710 9512
rect 22741 9503 22799 9509
rect 22741 9469 22753 9503
rect 22787 9500 22799 9503
rect 23308 9500 23336 9531
rect 24136 9512 24164 9540
rect 22787 9472 23336 9500
rect 23661 9503 23719 9509
rect 22787 9469 22799 9472
rect 22741 9463 22799 9469
rect 23661 9469 23673 9503
rect 23707 9469 23719 9503
rect 23661 9463 23719 9469
rect 21140 9404 22600 9432
rect 21140 9392 21146 9404
rect 18230 9364 18236 9376
rect 17972 9336 18236 9364
rect 18230 9324 18236 9336
rect 18288 9324 18294 9376
rect 19242 9324 19248 9376
rect 19300 9324 19306 9376
rect 19334 9324 19340 9376
rect 19392 9324 19398 9376
rect 20257 9367 20315 9373
rect 20257 9333 20269 9367
rect 20303 9364 20315 9367
rect 20806 9364 20812 9376
rect 20303 9336 20812 9364
rect 20303 9333 20315 9336
rect 20257 9327 20315 9333
rect 20806 9324 20812 9336
rect 20864 9324 20870 9376
rect 20990 9324 20996 9376
rect 21048 9364 21054 9376
rect 21174 9364 21180 9376
rect 21048 9336 21180 9364
rect 21048 9324 21054 9336
rect 21174 9324 21180 9336
rect 21232 9324 21238 9376
rect 22278 9324 22284 9376
rect 22336 9364 22342 9376
rect 22756 9364 22784 9463
rect 23382 9392 23388 9444
rect 23440 9432 23446 9444
rect 23676 9432 23704 9463
rect 24118 9460 24124 9512
rect 24176 9460 24182 9512
rect 23440 9404 23704 9432
rect 23440 9392 23446 9404
rect 22336 9336 22784 9364
rect 22336 9324 22342 9336
rect 1104 9274 28888 9296
rect 1104 9222 4423 9274
rect 4475 9222 4487 9274
rect 4539 9222 4551 9274
rect 4603 9222 4615 9274
rect 4667 9222 4679 9274
rect 4731 9222 11369 9274
rect 11421 9222 11433 9274
rect 11485 9222 11497 9274
rect 11549 9222 11561 9274
rect 11613 9222 11625 9274
rect 11677 9222 18315 9274
rect 18367 9222 18379 9274
rect 18431 9222 18443 9274
rect 18495 9222 18507 9274
rect 18559 9222 18571 9274
rect 18623 9222 25261 9274
rect 25313 9222 25325 9274
rect 25377 9222 25389 9274
rect 25441 9222 25453 9274
rect 25505 9222 25517 9274
rect 25569 9222 28888 9274
rect 1104 9200 28888 9222
rect 17770 9160 17776 9172
rect 15856 9132 17776 9160
rect 14369 9095 14427 9101
rect 14369 9061 14381 9095
rect 14415 9061 14427 9095
rect 14369 9055 14427 9061
rect 6886 8996 12434 9024
rect 934 8916 940 8968
rect 992 8956 998 8968
rect 1397 8959 1455 8965
rect 1397 8956 1409 8959
rect 992 8928 1409 8956
rect 992 8916 998 8928
rect 1397 8925 1409 8928
rect 1443 8925 1455 8959
rect 1397 8919 1455 8925
rect 1581 8823 1639 8829
rect 1581 8789 1593 8823
rect 1627 8820 1639 8823
rect 6886 8820 6914 8996
rect 12406 8888 12434 8996
rect 14277 8959 14335 8965
rect 14277 8925 14289 8959
rect 14323 8956 14335 8959
rect 14384 8956 14412 9055
rect 15010 8984 15016 9036
rect 15068 9024 15074 9036
rect 15856 9024 15884 9132
rect 17770 9120 17776 9132
rect 17828 9120 17834 9172
rect 18325 9163 18383 9169
rect 18325 9129 18337 9163
rect 18371 9160 18383 9163
rect 19242 9160 19248 9172
rect 18371 9132 19248 9160
rect 18371 9129 18383 9132
rect 18325 9123 18383 9129
rect 19242 9120 19248 9132
rect 19300 9120 19306 9172
rect 20254 9120 20260 9172
rect 20312 9160 20318 9172
rect 20441 9163 20499 9169
rect 20441 9160 20453 9163
rect 20312 9132 20453 9160
rect 20312 9120 20318 9132
rect 20441 9129 20453 9132
rect 20487 9129 20499 9163
rect 20441 9123 20499 9129
rect 20714 9120 20720 9172
rect 20772 9160 20778 9172
rect 20901 9163 20959 9169
rect 20901 9160 20913 9163
rect 20772 9132 20913 9160
rect 20772 9120 20778 9132
rect 20901 9129 20913 9132
rect 20947 9129 20959 9163
rect 20901 9123 20959 9129
rect 21085 9163 21143 9169
rect 21085 9129 21097 9163
rect 21131 9160 21143 9163
rect 21266 9160 21272 9172
rect 21131 9132 21272 9160
rect 21131 9129 21143 9132
rect 21085 9123 21143 9129
rect 21266 9120 21272 9132
rect 21324 9120 21330 9172
rect 22097 9163 22155 9169
rect 22097 9129 22109 9163
rect 22143 9129 22155 9163
rect 22097 9123 22155 9129
rect 17034 9052 17040 9104
rect 17092 9092 17098 9104
rect 19426 9092 19432 9104
rect 17092 9064 17264 9092
rect 17092 9052 17098 9064
rect 15068 8996 15884 9024
rect 15068 8984 15074 8996
rect 15930 8984 15936 9036
rect 15988 9024 15994 9036
rect 16485 9027 16543 9033
rect 16485 9024 16497 9027
rect 15988 8996 16497 9024
rect 15988 8984 15994 8996
rect 16485 8993 16497 8996
rect 16531 8993 16543 9027
rect 16485 8987 16543 8993
rect 17126 8984 17132 9036
rect 17184 8984 17190 9036
rect 17236 9024 17264 9064
rect 18432 9064 19432 9092
rect 17405 9027 17463 9033
rect 17405 9024 17417 9027
rect 17236 8996 17417 9024
rect 17405 8993 17417 8996
rect 17451 8993 17463 9027
rect 17405 8987 17463 8993
rect 17494 8984 17500 9036
rect 17552 9033 17558 9036
rect 17552 9027 17580 9033
rect 17568 8993 17580 9027
rect 17552 8987 17580 8993
rect 17552 8984 17558 8987
rect 17678 8984 17684 9036
rect 17736 9024 17742 9036
rect 18432 9024 18460 9064
rect 19426 9052 19432 9064
rect 19484 9052 19490 9104
rect 20806 9052 20812 9104
rect 20864 9092 20870 9104
rect 22002 9092 22008 9104
rect 20864 9064 22008 9092
rect 20864 9052 20870 9064
rect 22002 9052 22008 9064
rect 22060 9092 22066 9104
rect 22112 9092 22140 9123
rect 22278 9120 22284 9172
rect 22336 9120 22342 9172
rect 22060 9064 22140 9092
rect 23017 9095 23075 9101
rect 22060 9052 22066 9064
rect 23017 9061 23029 9095
rect 23063 9061 23075 9095
rect 23017 9055 23075 9061
rect 17736 8996 18460 9024
rect 17736 8984 17742 8996
rect 14323 8928 14412 8956
rect 14323 8925 14335 8928
rect 14277 8919 14335 8925
rect 16022 8916 16028 8968
rect 16080 8916 16086 8968
rect 16390 8916 16396 8968
rect 16448 8956 16454 8968
rect 18432 8965 18460 8996
rect 18874 8984 18880 9036
rect 18932 9024 18938 9036
rect 20717 9027 20775 9033
rect 18932 8996 20116 9024
rect 18932 8984 18938 8996
rect 16669 8959 16727 8965
rect 16669 8956 16681 8959
rect 16448 8928 16681 8956
rect 16448 8916 16454 8928
rect 16669 8925 16681 8928
rect 16715 8925 16727 8959
rect 16669 8919 16727 8925
rect 18417 8959 18475 8965
rect 18417 8925 18429 8959
rect 18463 8925 18475 8959
rect 18417 8919 18475 8925
rect 18598 8916 18604 8968
rect 18656 8916 18662 8968
rect 20088 8965 20116 8996
rect 20717 8993 20729 9027
rect 20763 9024 20775 9027
rect 20898 9024 20904 9036
rect 20763 8996 20904 9024
rect 20763 8993 20775 8996
rect 20717 8987 20775 8993
rect 20898 8984 20904 8996
rect 20956 9024 20962 9036
rect 21637 9027 21695 9033
rect 20956 8996 21128 9024
rect 20956 8984 20962 8996
rect 19337 8959 19395 8965
rect 19337 8925 19349 8959
rect 19383 8925 19395 8959
rect 19337 8919 19395 8925
rect 20073 8959 20131 8965
rect 20073 8925 20085 8959
rect 20119 8925 20131 8959
rect 20073 8919 20131 8925
rect 14734 8888 14740 8900
rect 12406 8860 14740 8888
rect 14734 8848 14740 8860
rect 14792 8848 14798 8900
rect 19352 8888 19380 8919
rect 20990 8916 20996 8968
rect 21048 8916 21054 8968
rect 21100 8956 21128 8996
rect 21637 8993 21649 9027
rect 21683 8993 21695 9027
rect 23032 9024 23060 9055
rect 23032 8996 23612 9024
rect 21637 8987 21695 8993
rect 21358 8956 21364 8968
rect 21100 8928 21364 8956
rect 21358 8916 21364 8928
rect 21416 8916 21422 8968
rect 21450 8916 21456 8968
rect 21508 8916 21514 8968
rect 20257 8891 20315 8897
rect 20257 8888 20269 8891
rect 19352 8860 20269 8888
rect 19352 8832 19380 8860
rect 20257 8857 20269 8860
rect 20303 8857 20315 8891
rect 21652 8888 21680 8987
rect 21818 8916 21824 8968
rect 21876 8956 21882 8968
rect 22373 8959 22431 8965
rect 22373 8956 22385 8959
rect 21876 8928 22385 8956
rect 21876 8916 21882 8928
rect 22373 8925 22385 8928
rect 22419 8956 22431 8959
rect 22646 8956 22652 8968
rect 22419 8928 22652 8956
rect 22419 8925 22431 8928
rect 22373 8919 22431 8925
rect 22646 8916 22652 8928
rect 22704 8916 22710 8968
rect 23109 8959 23167 8965
rect 23109 8925 23121 8959
rect 23155 8925 23167 8959
rect 23109 8919 23167 8925
rect 23293 8959 23351 8965
rect 23293 8925 23305 8959
rect 23339 8956 23351 8959
rect 23382 8956 23388 8968
rect 23339 8928 23388 8956
rect 23339 8925 23351 8928
rect 23293 8919 23351 8925
rect 20257 8851 20315 8857
rect 21468 8860 21680 8888
rect 21913 8891 21971 8897
rect 21468 8832 21496 8860
rect 21913 8857 21925 8891
rect 21959 8857 21971 8891
rect 21913 8851 21971 8857
rect 22129 8891 22187 8897
rect 22129 8857 22141 8891
rect 22175 8888 22187 8891
rect 22175 8860 22784 8888
rect 22175 8857 22187 8860
rect 22129 8851 22187 8857
rect 1627 8792 6914 8820
rect 1627 8789 1639 8792
rect 1581 8783 1639 8789
rect 14090 8780 14096 8832
rect 14148 8780 14154 8832
rect 14829 8823 14887 8829
rect 14829 8789 14841 8823
rect 14875 8820 14887 8823
rect 15289 8823 15347 8829
rect 15289 8820 15301 8823
rect 14875 8792 15301 8820
rect 14875 8789 14887 8792
rect 14829 8783 14887 8789
rect 15289 8789 15301 8792
rect 15335 8789 15347 8823
rect 15289 8783 15347 8789
rect 16206 8780 16212 8832
rect 16264 8780 16270 8832
rect 18230 8780 18236 8832
rect 18288 8820 18294 8832
rect 18417 8823 18475 8829
rect 18417 8820 18429 8823
rect 18288 8792 18429 8820
rect 18288 8780 18294 8792
rect 18417 8789 18429 8792
rect 18463 8789 18475 8823
rect 18417 8783 18475 8789
rect 19334 8780 19340 8832
rect 19392 8780 19398 8832
rect 19981 8823 20039 8829
rect 19981 8789 19993 8823
rect 20027 8820 20039 8823
rect 20346 8820 20352 8832
rect 20027 8792 20352 8820
rect 20027 8789 20039 8792
rect 19981 8783 20039 8789
rect 20346 8780 20352 8792
rect 20404 8780 20410 8832
rect 20530 8780 20536 8832
rect 20588 8820 20594 8832
rect 20717 8823 20775 8829
rect 20717 8820 20729 8823
rect 20588 8792 20729 8820
rect 20588 8780 20594 8792
rect 20717 8789 20729 8792
rect 20763 8789 20775 8823
rect 20717 8783 20775 8789
rect 21450 8780 21456 8832
rect 21508 8780 21514 8832
rect 21542 8780 21548 8832
rect 21600 8780 21606 8832
rect 21928 8820 21956 8851
rect 22462 8820 22468 8832
rect 21928 8792 22468 8820
rect 22462 8780 22468 8792
rect 22520 8780 22526 8832
rect 22646 8780 22652 8832
rect 22704 8780 22710 8832
rect 22756 8829 22784 8860
rect 22830 8848 22836 8900
rect 22888 8897 22894 8900
rect 22888 8891 22916 8897
rect 22904 8888 22916 8891
rect 23124 8888 23152 8919
rect 23382 8916 23388 8928
rect 23440 8916 23446 8968
rect 23584 8965 23612 8996
rect 23569 8959 23627 8965
rect 23569 8925 23581 8959
rect 23615 8925 23627 8959
rect 23569 8919 23627 8925
rect 24673 8959 24731 8965
rect 24673 8925 24685 8959
rect 24719 8956 24731 8959
rect 24762 8956 24768 8968
rect 24719 8928 24768 8956
rect 24719 8925 24731 8928
rect 24673 8919 24731 8925
rect 24762 8916 24768 8928
rect 24820 8916 24826 8968
rect 22904 8860 24164 8888
rect 22904 8857 22916 8860
rect 22888 8851 22916 8857
rect 22888 8848 22894 8851
rect 24136 8832 24164 8860
rect 22741 8823 22799 8829
rect 22741 8789 22753 8823
rect 22787 8820 22799 8823
rect 23474 8820 23480 8832
rect 22787 8792 23480 8820
rect 22787 8789 22799 8792
rect 22741 8783 22799 8789
rect 23474 8780 23480 8792
rect 23532 8780 23538 8832
rect 23750 8780 23756 8832
rect 23808 8780 23814 8832
rect 24118 8780 24124 8832
rect 24176 8820 24182 8832
rect 24489 8823 24547 8829
rect 24489 8820 24501 8823
rect 24176 8792 24501 8820
rect 24176 8780 24182 8792
rect 24489 8789 24501 8792
rect 24535 8789 24547 8823
rect 24489 8783 24547 8789
rect 1104 8730 28888 8752
rect 1104 8678 5083 8730
rect 5135 8678 5147 8730
rect 5199 8678 5211 8730
rect 5263 8678 5275 8730
rect 5327 8678 5339 8730
rect 5391 8678 12029 8730
rect 12081 8678 12093 8730
rect 12145 8678 12157 8730
rect 12209 8678 12221 8730
rect 12273 8678 12285 8730
rect 12337 8678 18975 8730
rect 19027 8678 19039 8730
rect 19091 8678 19103 8730
rect 19155 8678 19167 8730
rect 19219 8678 19231 8730
rect 19283 8678 25921 8730
rect 25973 8678 25985 8730
rect 26037 8678 26049 8730
rect 26101 8678 26113 8730
rect 26165 8678 26177 8730
rect 26229 8678 28888 8730
rect 1104 8656 28888 8678
rect 15102 8616 15108 8628
rect 13924 8588 15108 8616
rect 13924 8489 13952 8588
rect 15102 8576 15108 8588
rect 15160 8576 15166 8628
rect 15657 8619 15715 8625
rect 15657 8585 15669 8619
rect 15703 8616 15715 8619
rect 15930 8616 15936 8628
rect 15703 8588 15936 8616
rect 15703 8585 15715 8588
rect 15657 8579 15715 8585
rect 15930 8576 15936 8588
rect 15988 8576 15994 8628
rect 16022 8576 16028 8628
rect 16080 8616 16086 8628
rect 16669 8619 16727 8625
rect 16669 8616 16681 8619
rect 16080 8588 16681 8616
rect 16080 8576 16086 8588
rect 16669 8585 16681 8588
rect 16715 8585 16727 8619
rect 18233 8619 18291 8625
rect 16669 8579 16727 8585
rect 16960 8588 18184 8616
rect 14090 8508 14096 8560
rect 14148 8548 14154 8560
rect 14185 8551 14243 8557
rect 14185 8548 14197 8551
rect 14148 8520 14197 8548
rect 14148 8508 14154 8520
rect 14185 8517 14197 8520
rect 14231 8517 14243 8551
rect 15746 8548 15752 8560
rect 15410 8520 15752 8548
rect 14185 8511 14243 8517
rect 15746 8508 15752 8520
rect 15804 8508 15810 8560
rect 16301 8551 16359 8557
rect 16301 8517 16313 8551
rect 16347 8548 16359 8551
rect 16960 8548 16988 8588
rect 18156 8560 18184 8588
rect 18233 8585 18245 8619
rect 18279 8616 18291 8619
rect 19334 8616 19340 8628
rect 18279 8588 19340 8616
rect 18279 8585 18291 8588
rect 18233 8579 18291 8585
rect 19334 8576 19340 8588
rect 19392 8576 19398 8628
rect 20346 8576 20352 8628
rect 20404 8576 20410 8628
rect 20806 8576 20812 8628
rect 20864 8576 20870 8628
rect 21361 8619 21419 8625
rect 21361 8585 21373 8619
rect 21407 8616 21419 8619
rect 21407 8588 21496 8616
rect 21407 8585 21419 8588
rect 21361 8579 21419 8585
rect 16347 8520 16988 8548
rect 17037 8551 17095 8557
rect 16347 8517 16359 8520
rect 16301 8511 16359 8517
rect 17037 8517 17049 8551
rect 17083 8548 17095 8551
rect 17218 8548 17224 8560
rect 17083 8520 17224 8548
rect 17083 8517 17095 8520
rect 17037 8511 17095 8517
rect 17218 8508 17224 8520
rect 17276 8508 17282 8560
rect 18138 8508 18144 8560
rect 18196 8508 18202 8560
rect 18690 8508 18696 8560
rect 18748 8508 18754 8560
rect 13909 8483 13967 8489
rect 13909 8449 13921 8483
rect 13955 8449 13967 8483
rect 15764 8480 15792 8508
rect 15933 8483 15991 8489
rect 15933 8480 15945 8483
rect 15764 8452 15945 8480
rect 13909 8443 13967 8449
rect 15933 8449 15945 8452
rect 15979 8449 15991 8483
rect 15933 8443 15991 8449
rect 17129 8483 17187 8489
rect 17129 8449 17141 8483
rect 17175 8480 17187 8483
rect 17497 8483 17555 8489
rect 17497 8480 17509 8483
rect 17175 8452 17509 8480
rect 17175 8449 17187 8452
rect 17129 8443 17187 8449
rect 17497 8449 17509 8452
rect 17543 8449 17555 8483
rect 17770 8480 17776 8492
rect 17497 8443 17555 8449
rect 17604 8452 17776 8480
rect 16390 8372 16396 8424
rect 16448 8372 16454 8424
rect 17313 8415 17371 8421
rect 17313 8381 17325 8415
rect 17359 8412 17371 8415
rect 17604 8412 17632 8452
rect 17770 8440 17776 8452
rect 17828 8480 17834 8492
rect 17828 8452 18184 8480
rect 17828 8440 17834 8452
rect 17359 8384 17632 8412
rect 18049 8415 18107 8421
rect 17359 8381 17371 8384
rect 17313 8375 17371 8381
rect 18049 8381 18061 8415
rect 18095 8381 18107 8415
rect 18049 8375 18107 8381
rect 16408 8344 16436 8372
rect 18064 8344 18092 8375
rect 16408 8316 18092 8344
rect 18156 8276 18184 8452
rect 19978 8440 19984 8492
rect 20036 8440 20042 8492
rect 20254 8440 20260 8492
rect 20312 8440 20318 8492
rect 20364 8489 20392 8576
rect 20824 8548 20852 8576
rect 20824 8520 20944 8548
rect 20916 8489 20944 8520
rect 21468 8492 21496 8588
rect 21542 8576 21548 8628
rect 21600 8576 21606 8628
rect 22002 8576 22008 8628
rect 22060 8616 22066 8628
rect 22060 8576 22094 8616
rect 22646 8576 22652 8628
rect 22704 8616 22710 8628
rect 22833 8619 22891 8625
rect 22833 8616 22845 8619
rect 22704 8588 22845 8616
rect 22704 8576 22710 8588
rect 22833 8585 22845 8588
rect 22879 8585 22891 8619
rect 22833 8579 22891 8585
rect 23201 8619 23259 8625
rect 23201 8585 23213 8619
rect 23247 8616 23259 8619
rect 23382 8616 23388 8628
rect 23247 8588 23388 8616
rect 23247 8585 23259 8588
rect 23201 8579 23259 8585
rect 23382 8576 23388 8588
rect 23440 8576 23446 8628
rect 23750 8616 23756 8628
rect 23584 8588 23756 8616
rect 21560 8548 21588 8576
rect 22066 8548 22094 8576
rect 22925 8551 22983 8557
rect 22925 8548 22937 8551
rect 21560 8520 21956 8548
rect 22066 8520 22937 8548
rect 20349 8483 20407 8489
rect 20349 8449 20361 8483
rect 20395 8449 20407 8483
rect 20349 8443 20407 8449
rect 20625 8483 20683 8489
rect 20625 8449 20637 8483
rect 20671 8480 20683 8483
rect 20809 8483 20867 8489
rect 20809 8480 20821 8483
rect 20671 8452 20821 8480
rect 20671 8449 20683 8452
rect 20625 8443 20683 8449
rect 20809 8449 20821 8452
rect 20855 8449 20867 8483
rect 20809 8443 20867 8449
rect 20901 8483 20959 8489
rect 20901 8449 20913 8483
rect 20947 8449 20959 8483
rect 20901 8443 20959 8449
rect 21082 8440 21088 8492
rect 21140 8480 21146 8492
rect 21269 8483 21327 8489
rect 21269 8480 21281 8483
rect 21140 8452 21281 8480
rect 21140 8440 21146 8452
rect 21269 8449 21281 8452
rect 21315 8449 21327 8483
rect 21269 8443 21327 8449
rect 21450 8440 21456 8492
rect 21508 8480 21514 8492
rect 21508 8452 21606 8480
rect 21508 8440 21514 8452
rect 19705 8415 19763 8421
rect 19705 8381 19717 8415
rect 19751 8412 19763 8415
rect 20073 8415 20131 8421
rect 20073 8412 20085 8415
rect 19751 8384 20085 8412
rect 19751 8381 19763 8384
rect 19705 8375 19763 8381
rect 20073 8381 20085 8384
rect 20119 8381 20131 8415
rect 20073 8375 20131 8381
rect 20162 8372 20168 8424
rect 20220 8412 20226 8424
rect 20530 8412 20536 8424
rect 20220 8384 20536 8412
rect 20220 8372 20226 8384
rect 20530 8372 20536 8384
rect 20588 8372 20594 8424
rect 21174 8372 21180 8424
rect 21232 8372 21238 8424
rect 21578 8412 21606 8452
rect 21634 8440 21640 8492
rect 21692 8440 21698 8492
rect 21821 8483 21879 8489
rect 21821 8449 21833 8483
rect 21867 8449 21879 8483
rect 21928 8480 21956 8520
rect 22925 8517 22937 8520
rect 22971 8517 22983 8551
rect 22925 8511 22983 8517
rect 23017 8551 23075 8557
rect 23017 8517 23029 8551
rect 23063 8548 23075 8551
rect 23474 8548 23480 8560
rect 23063 8520 23480 8548
rect 23063 8517 23075 8520
rect 23017 8511 23075 8517
rect 23474 8508 23480 8520
rect 23532 8508 23538 8560
rect 23584 8557 23612 8588
rect 23750 8576 23756 8588
rect 23808 8576 23814 8628
rect 23569 8551 23627 8557
rect 23569 8517 23581 8551
rect 23615 8517 23627 8551
rect 23569 8511 23627 8517
rect 24026 8508 24032 8560
rect 24084 8508 24090 8560
rect 22465 8483 22523 8489
rect 22465 8480 22477 8483
rect 21928 8452 22477 8480
rect 21821 8443 21879 8449
rect 22465 8449 22477 8452
rect 22511 8449 22523 8483
rect 22465 8443 22523 8449
rect 21836 8412 21864 8443
rect 21284 8384 21496 8412
rect 21578 8384 21864 8412
rect 22480 8412 22508 8443
rect 22554 8440 22560 8492
rect 22612 8480 22618 8492
rect 22649 8483 22707 8489
rect 22649 8480 22661 8483
rect 22612 8452 22661 8480
rect 22612 8440 22618 8452
rect 22649 8449 22661 8452
rect 22695 8449 22707 8483
rect 22649 8443 22707 8449
rect 22480 8384 22692 8412
rect 21284 8276 21312 8384
rect 21468 8344 21496 8384
rect 21913 8347 21971 8353
rect 21913 8344 21925 8347
rect 21468 8316 21925 8344
rect 21913 8313 21925 8316
rect 21959 8313 21971 8347
rect 22664 8344 22692 8384
rect 23198 8372 23204 8424
rect 23256 8412 23262 8424
rect 23293 8415 23351 8421
rect 23293 8412 23305 8415
rect 23256 8384 23305 8412
rect 23256 8372 23262 8384
rect 23293 8381 23305 8384
rect 23339 8381 23351 8415
rect 23293 8375 23351 8381
rect 25041 8347 25099 8353
rect 25041 8344 25053 8347
rect 22664 8316 23428 8344
rect 21913 8307 21971 8313
rect 18156 8248 21312 8276
rect 23400 8276 23428 8316
rect 24780 8316 25053 8344
rect 24780 8288 24808 8316
rect 25041 8313 25053 8316
rect 25087 8313 25099 8347
rect 25041 8307 25099 8313
rect 24210 8276 24216 8288
rect 23400 8248 24216 8276
rect 24210 8236 24216 8248
rect 24268 8236 24274 8288
rect 24762 8236 24768 8288
rect 24820 8236 24826 8288
rect 1104 8186 28888 8208
rect 1104 8134 4423 8186
rect 4475 8134 4487 8186
rect 4539 8134 4551 8186
rect 4603 8134 4615 8186
rect 4667 8134 4679 8186
rect 4731 8134 11369 8186
rect 11421 8134 11433 8186
rect 11485 8134 11497 8186
rect 11549 8134 11561 8186
rect 11613 8134 11625 8186
rect 11677 8134 18315 8186
rect 18367 8134 18379 8186
rect 18431 8134 18443 8186
rect 18495 8134 18507 8186
rect 18559 8134 18571 8186
rect 18623 8134 25261 8186
rect 25313 8134 25325 8186
rect 25377 8134 25389 8186
rect 25441 8134 25453 8186
rect 25505 8134 25517 8186
rect 25569 8134 28888 8186
rect 1104 8112 28888 8134
rect 15102 8032 15108 8084
rect 15160 8072 15166 8084
rect 15933 8075 15991 8081
rect 15933 8072 15945 8075
rect 15160 8044 15945 8072
rect 15160 8032 15166 8044
rect 15933 8041 15945 8044
rect 15979 8041 15991 8075
rect 15933 8035 15991 8041
rect 17126 8032 17132 8084
rect 17184 8072 17190 8084
rect 17494 8072 17500 8084
rect 17184 8044 17500 8072
rect 17184 8032 17190 8044
rect 17494 8032 17500 8044
rect 17552 8072 17558 8084
rect 18690 8072 18696 8084
rect 17552 8044 18696 8072
rect 17552 8032 17558 8044
rect 18690 8032 18696 8044
rect 18748 8072 18754 8084
rect 19245 8075 19303 8081
rect 18748 8044 19012 8072
rect 18748 8032 18754 8044
rect 17862 8004 17868 8016
rect 17420 7976 17868 8004
rect 17420 7877 17448 7976
rect 17862 7964 17868 7976
rect 17920 7964 17926 8016
rect 18322 8004 18328 8016
rect 18248 7976 18328 8004
rect 18141 7939 18199 7945
rect 18141 7905 18153 7939
rect 18187 7936 18199 7939
rect 18248 7936 18276 7976
rect 18322 7964 18328 7976
rect 18380 7964 18386 8016
rect 18984 7945 19012 8044
rect 19245 8041 19257 8075
rect 19291 8072 19303 8075
rect 20254 8072 20260 8084
rect 19291 8044 20260 8072
rect 19291 8041 19303 8044
rect 19245 8035 19303 8041
rect 20254 8032 20260 8044
rect 20312 8032 20318 8084
rect 20533 8075 20591 8081
rect 20533 8041 20545 8075
rect 20579 8072 20591 8075
rect 20579 8044 20852 8072
rect 20579 8041 20591 8044
rect 20533 8035 20591 8041
rect 20824 8016 20852 8044
rect 21174 8032 21180 8084
rect 21232 8072 21238 8084
rect 22830 8072 22836 8084
rect 21232 8044 22836 8072
rect 21232 8032 21238 8044
rect 22830 8032 22836 8044
rect 22888 8032 22894 8084
rect 23474 8032 23480 8084
rect 23532 8072 23538 8084
rect 23753 8075 23811 8081
rect 23753 8072 23765 8075
rect 23532 8044 23765 8072
rect 23532 8032 23538 8044
rect 23753 8041 23765 8044
rect 23799 8041 23811 8075
rect 23753 8035 23811 8041
rect 23934 8032 23940 8084
rect 23992 8032 23998 8084
rect 24489 8075 24547 8081
rect 24489 8041 24501 8075
rect 24535 8072 24547 8075
rect 24762 8072 24768 8084
rect 24535 8044 24768 8072
rect 24535 8041 24547 8044
rect 24489 8035 24547 8041
rect 24762 8032 24768 8044
rect 24820 8032 24826 8084
rect 19889 8007 19947 8013
rect 19889 7973 19901 8007
rect 19935 8004 19947 8007
rect 20714 8004 20720 8016
rect 19935 7976 20720 8004
rect 19935 7973 19947 7976
rect 19889 7967 19947 7973
rect 20714 7964 20720 7976
rect 20772 7964 20778 8016
rect 20806 7964 20812 8016
rect 20864 8004 20870 8016
rect 20864 7976 21956 8004
rect 20864 7964 20870 7976
rect 18187 7908 18276 7936
rect 18969 7939 19027 7945
rect 18187 7905 18199 7908
rect 18141 7899 18199 7905
rect 18969 7905 18981 7939
rect 19015 7936 19027 7939
rect 19981 7939 20039 7945
rect 19015 7908 19656 7936
rect 19015 7905 19027 7908
rect 18969 7899 19027 7905
rect 17405 7871 17463 7877
rect 17405 7837 17417 7871
rect 17451 7837 17463 7871
rect 17405 7831 17463 7837
rect 17678 7828 17684 7880
rect 17736 7828 17742 7880
rect 17770 7828 17776 7880
rect 17828 7828 17834 7880
rect 17865 7871 17923 7877
rect 17865 7837 17877 7871
rect 17911 7868 17923 7871
rect 18230 7868 18236 7880
rect 17911 7840 18236 7868
rect 17911 7837 17923 7840
rect 17865 7831 17923 7837
rect 18230 7828 18236 7840
rect 18288 7828 18294 7880
rect 18690 7828 18696 7880
rect 18748 7828 18754 7880
rect 19426 7828 19432 7880
rect 19484 7868 19490 7880
rect 19628 7877 19656 7908
rect 19981 7905 19993 7939
rect 20027 7936 20039 7939
rect 20990 7936 20996 7948
rect 20027 7908 20996 7936
rect 20027 7905 20039 7908
rect 19981 7899 20039 7905
rect 20990 7896 20996 7908
rect 21048 7896 21054 7948
rect 19521 7871 19579 7877
rect 19521 7868 19533 7871
rect 19484 7840 19533 7868
rect 19484 7828 19490 7840
rect 19521 7837 19533 7840
rect 19567 7837 19579 7871
rect 19521 7831 19579 7837
rect 19613 7871 19671 7877
rect 19613 7837 19625 7871
rect 19659 7868 19671 7871
rect 20070 7868 20076 7880
rect 19659 7840 20076 7868
rect 19659 7837 19671 7840
rect 19613 7831 19671 7837
rect 20070 7828 20076 7840
rect 20128 7868 20134 7880
rect 20898 7868 20904 7880
rect 20128 7840 20484 7868
rect 20128 7828 20134 7840
rect 20456 7812 20484 7840
rect 20548 7840 20904 7868
rect 18003 7803 18061 7809
rect 18003 7769 18015 7803
rect 18049 7800 18061 7803
rect 18785 7803 18843 7809
rect 18785 7800 18797 7803
rect 18049 7772 18797 7800
rect 18049 7769 18061 7772
rect 18003 7763 18061 7769
rect 18785 7769 18797 7772
rect 18831 7800 18843 7803
rect 20162 7800 20168 7812
rect 18831 7772 20168 7800
rect 18831 7769 18843 7772
rect 18785 7763 18843 7769
rect 20162 7760 20168 7772
rect 20220 7760 20226 7812
rect 20438 7760 20444 7812
rect 20496 7760 20502 7812
rect 17034 7692 17040 7744
rect 17092 7732 17098 7744
rect 17497 7735 17555 7741
rect 17497 7732 17509 7735
rect 17092 7704 17509 7732
rect 17092 7692 17098 7704
rect 17497 7701 17509 7704
rect 17543 7701 17555 7735
rect 17497 7695 17555 7701
rect 18230 7692 18236 7744
rect 18288 7732 18294 7744
rect 18325 7735 18383 7741
rect 18325 7732 18337 7735
rect 18288 7704 18337 7732
rect 18288 7692 18294 7704
rect 18325 7701 18337 7704
rect 18371 7701 18383 7735
rect 18325 7695 18383 7701
rect 19705 7735 19763 7741
rect 19705 7701 19717 7735
rect 19751 7732 19763 7735
rect 20548 7732 20576 7840
rect 20898 7828 20904 7840
rect 20956 7828 20962 7880
rect 21818 7828 21824 7880
rect 21876 7828 21882 7880
rect 21928 7809 21956 7976
rect 22462 7964 22468 8016
rect 22520 8004 22526 8016
rect 22520 7976 24992 8004
rect 22520 7964 22526 7976
rect 24026 7896 24032 7948
rect 24084 7896 24090 7948
rect 24118 7896 24124 7948
rect 24176 7896 24182 7948
rect 24504 7908 24808 7936
rect 23937 7871 23995 7877
rect 23937 7837 23949 7871
rect 23983 7837 23995 7871
rect 24044 7868 24072 7896
rect 24397 7871 24455 7877
rect 24397 7868 24409 7871
rect 24044 7840 24409 7868
rect 23937 7831 23995 7837
rect 24397 7837 24409 7840
rect 24443 7837 24455 7871
rect 24397 7831 24455 7837
rect 21913 7803 21971 7809
rect 21913 7769 21925 7803
rect 21959 7769 21971 7803
rect 21913 7763 21971 7769
rect 19751 7704 20576 7732
rect 19751 7701 19763 7704
rect 19705 7695 19763 7701
rect 20714 7692 20720 7744
rect 20772 7732 20778 7744
rect 22554 7732 22560 7744
rect 20772 7704 22560 7732
rect 20772 7692 20778 7704
rect 22554 7692 22560 7704
rect 22612 7692 22618 7744
rect 23198 7692 23204 7744
rect 23256 7692 23262 7744
rect 23952 7732 23980 7831
rect 24210 7760 24216 7812
rect 24268 7800 24274 7812
rect 24504 7800 24532 7908
rect 24673 7871 24731 7877
rect 24673 7837 24685 7871
rect 24719 7837 24731 7871
rect 24673 7831 24731 7837
rect 24268 7772 24532 7800
rect 24268 7760 24274 7772
rect 24302 7732 24308 7744
rect 23952 7704 24308 7732
rect 24302 7692 24308 7704
rect 24360 7732 24366 7744
rect 24688 7732 24716 7831
rect 24780 7800 24808 7908
rect 24964 7877 24992 7976
rect 24949 7871 25007 7877
rect 24949 7837 24961 7871
rect 24995 7837 25007 7871
rect 24949 7831 25007 7837
rect 28258 7800 28264 7812
rect 24780 7772 28264 7800
rect 28258 7760 28264 7772
rect 28316 7760 28322 7812
rect 24360 7704 24716 7732
rect 24360 7692 24366 7704
rect 24854 7692 24860 7744
rect 24912 7692 24918 7744
rect 25038 7692 25044 7744
rect 25096 7732 25102 7744
rect 25133 7735 25191 7741
rect 25133 7732 25145 7735
rect 25096 7704 25145 7732
rect 25096 7692 25102 7704
rect 25133 7701 25145 7704
rect 25179 7701 25191 7735
rect 25133 7695 25191 7701
rect 1104 7642 28888 7664
rect 1104 7590 5083 7642
rect 5135 7590 5147 7642
rect 5199 7590 5211 7642
rect 5263 7590 5275 7642
rect 5327 7590 5339 7642
rect 5391 7590 12029 7642
rect 12081 7590 12093 7642
rect 12145 7590 12157 7642
rect 12209 7590 12221 7642
rect 12273 7590 12285 7642
rect 12337 7590 18975 7642
rect 19027 7590 19039 7642
rect 19091 7590 19103 7642
rect 19155 7590 19167 7642
rect 19219 7590 19231 7642
rect 19283 7590 25921 7642
rect 25973 7590 25985 7642
rect 26037 7590 26049 7642
rect 26101 7590 26113 7642
rect 26165 7590 26177 7642
rect 26229 7590 28888 7642
rect 1104 7568 28888 7590
rect 14737 7531 14795 7537
rect 14737 7497 14749 7531
rect 14783 7528 14795 7531
rect 16390 7528 16396 7540
rect 14783 7500 16396 7528
rect 14783 7497 14795 7500
rect 14737 7491 14795 7497
rect 16390 7488 16396 7500
rect 16448 7488 16454 7540
rect 17494 7528 17500 7540
rect 17236 7500 17500 7528
rect 15746 7420 15752 7472
rect 15804 7420 15810 7472
rect 16206 7420 16212 7472
rect 16264 7420 16270 7472
rect 17236 7469 17264 7500
rect 17494 7488 17500 7500
rect 17552 7488 17558 7540
rect 17589 7531 17647 7537
rect 17589 7497 17601 7531
rect 17635 7528 17647 7531
rect 17678 7528 17684 7540
rect 17635 7500 17684 7528
rect 17635 7497 17647 7500
rect 17589 7491 17647 7497
rect 17678 7488 17684 7500
rect 17736 7488 17742 7540
rect 18322 7488 18328 7540
rect 18380 7488 18386 7540
rect 18690 7488 18696 7540
rect 18748 7528 18754 7540
rect 20714 7537 20720 7540
rect 20533 7531 20591 7537
rect 20533 7528 20545 7531
rect 18748 7500 20545 7528
rect 18748 7488 18754 7500
rect 20533 7497 20545 7500
rect 20579 7497 20591 7531
rect 20533 7491 20591 7497
rect 20701 7531 20720 7537
rect 20701 7497 20713 7531
rect 20701 7491 20720 7497
rect 20714 7488 20720 7491
rect 20772 7488 20778 7540
rect 20990 7488 20996 7540
rect 21048 7528 21054 7540
rect 21085 7531 21143 7537
rect 21085 7528 21097 7531
rect 21048 7500 21097 7528
rect 21048 7488 21054 7500
rect 21085 7497 21097 7500
rect 21131 7497 21143 7531
rect 21085 7491 21143 7497
rect 22462 7488 22468 7540
rect 22520 7488 22526 7540
rect 17221 7463 17279 7469
rect 17221 7429 17233 7463
rect 17267 7429 17279 7463
rect 17221 7423 17279 7429
rect 17405 7463 17463 7469
rect 17405 7429 17417 7463
rect 17451 7429 17463 7463
rect 17405 7423 17463 7429
rect 17420 7392 17448 7423
rect 19702 7420 19708 7472
rect 19760 7420 19766 7472
rect 20438 7420 20444 7472
rect 20496 7420 20502 7472
rect 20901 7463 20959 7469
rect 20901 7429 20913 7463
rect 20947 7429 20959 7463
rect 20901 7423 20959 7429
rect 17586 7392 17592 7404
rect 17420 7364 17592 7392
rect 17586 7352 17592 7364
rect 17644 7392 17650 7404
rect 17681 7395 17739 7401
rect 17681 7392 17693 7395
rect 17644 7364 17693 7392
rect 17644 7352 17650 7364
rect 17681 7361 17693 7364
rect 17727 7361 17739 7395
rect 20916 7392 20944 7423
rect 21450 7420 21456 7472
rect 21508 7420 21514 7472
rect 21174 7392 21180 7404
rect 20916 7364 21180 7392
rect 17681 7355 17739 7361
rect 21174 7352 21180 7364
rect 21232 7352 21238 7404
rect 21634 7352 21640 7404
rect 21692 7352 21698 7404
rect 21821 7395 21879 7401
rect 21821 7361 21833 7395
rect 21867 7361 21879 7395
rect 21821 7355 21879 7361
rect 16485 7327 16543 7333
rect 16485 7293 16497 7327
rect 16531 7324 16543 7327
rect 16574 7324 16580 7336
rect 16531 7296 16580 7324
rect 16531 7293 16543 7296
rect 16485 7287 16543 7293
rect 16574 7284 16580 7296
rect 16632 7284 16638 7336
rect 18417 7327 18475 7333
rect 18417 7293 18429 7327
rect 18463 7293 18475 7327
rect 18417 7287 18475 7293
rect 16592 7256 16620 7284
rect 18432 7256 18460 7287
rect 18690 7284 18696 7336
rect 18748 7284 18754 7336
rect 21836 7324 21864 7355
rect 21910 7352 21916 7404
rect 21968 7352 21974 7404
rect 22097 7395 22155 7401
rect 22097 7361 22109 7395
rect 22143 7361 22155 7395
rect 22097 7355 22155 7361
rect 21284 7296 21864 7324
rect 22112 7324 22140 7355
rect 22186 7352 22192 7404
rect 22244 7352 22250 7404
rect 22281 7395 22339 7401
rect 22281 7361 22293 7395
rect 22327 7392 22339 7395
rect 22327 7364 22784 7392
rect 24794 7364 24900 7392
rect 22327 7361 22339 7364
rect 22281 7355 22339 7361
rect 22756 7336 22784 7364
rect 22370 7324 22376 7336
rect 22112 7296 22376 7324
rect 20898 7256 20904 7268
rect 16592 7228 18460 7256
rect 20732 7228 20904 7256
rect 20732 7197 20760 7228
rect 20898 7216 20904 7228
rect 20956 7216 20962 7268
rect 20717 7191 20775 7197
rect 20717 7157 20729 7191
rect 20763 7157 20775 7191
rect 20717 7151 20775 7157
rect 21174 7148 21180 7200
rect 21232 7188 21238 7200
rect 21284 7197 21312 7296
rect 22370 7284 22376 7296
rect 22428 7284 22434 7336
rect 22554 7284 22560 7336
rect 22612 7284 22618 7336
rect 22738 7284 22744 7336
rect 22796 7284 22802 7336
rect 22830 7284 22836 7336
rect 22888 7284 22894 7336
rect 22925 7327 22983 7333
rect 22925 7293 22937 7327
rect 22971 7293 22983 7327
rect 22925 7287 22983 7293
rect 22940 7256 22968 7287
rect 23014 7284 23020 7336
rect 23072 7284 23078 7336
rect 23198 7284 23204 7336
rect 23256 7324 23262 7336
rect 23385 7327 23443 7333
rect 23385 7324 23397 7327
rect 23256 7296 23397 7324
rect 23256 7284 23262 7296
rect 23385 7293 23397 7296
rect 23431 7293 23443 7327
rect 23385 7287 23443 7293
rect 23658 7284 23664 7336
rect 23716 7284 23722 7336
rect 24872 7268 24900 7364
rect 22572 7228 22968 7256
rect 22572 7200 22600 7228
rect 21269 7191 21327 7197
rect 21269 7188 21281 7191
rect 21232 7160 21281 7188
rect 21232 7148 21238 7160
rect 21269 7157 21281 7160
rect 21315 7157 21327 7191
rect 21269 7151 21327 7157
rect 22554 7148 22560 7200
rect 22612 7148 22618 7200
rect 22940 7188 22968 7228
rect 24854 7216 24860 7268
rect 24912 7216 24918 7268
rect 24946 7188 24952 7200
rect 22940 7160 24952 7188
rect 24946 7148 24952 7160
rect 25004 7188 25010 7200
rect 25133 7191 25191 7197
rect 25133 7188 25145 7191
rect 25004 7160 25145 7188
rect 25004 7148 25010 7160
rect 25133 7157 25145 7160
rect 25179 7157 25191 7191
rect 25133 7151 25191 7157
rect 1104 7098 28888 7120
rect 1104 7046 4423 7098
rect 4475 7046 4487 7098
rect 4539 7046 4551 7098
rect 4603 7046 4615 7098
rect 4667 7046 4679 7098
rect 4731 7046 11369 7098
rect 11421 7046 11433 7098
rect 11485 7046 11497 7098
rect 11549 7046 11561 7098
rect 11613 7046 11625 7098
rect 11677 7046 18315 7098
rect 18367 7046 18379 7098
rect 18431 7046 18443 7098
rect 18495 7046 18507 7098
rect 18559 7046 18571 7098
rect 18623 7046 25261 7098
rect 25313 7046 25325 7098
rect 25377 7046 25389 7098
rect 25441 7046 25453 7098
rect 25505 7046 25517 7098
rect 25569 7046 28888 7098
rect 1104 7024 28888 7046
rect 16656 6987 16714 6993
rect 16656 6953 16668 6987
rect 16702 6984 16714 6987
rect 17034 6984 17040 6996
rect 16702 6956 17040 6984
rect 16702 6953 16714 6956
rect 16656 6947 16714 6953
rect 17034 6944 17040 6956
rect 17092 6944 17098 6996
rect 17678 6944 17684 6996
rect 17736 6984 17742 6996
rect 18141 6987 18199 6993
rect 18141 6984 18153 6987
rect 17736 6956 18153 6984
rect 17736 6944 17742 6956
rect 18141 6953 18153 6956
rect 18187 6953 18199 6987
rect 18141 6947 18199 6953
rect 18690 6944 18696 6996
rect 18748 6944 18754 6996
rect 21563 6987 21621 6993
rect 21563 6953 21575 6987
rect 21609 6984 21621 6987
rect 23293 6987 23351 6993
rect 23293 6984 23305 6987
rect 21609 6956 23305 6984
rect 21609 6953 21621 6956
rect 21563 6947 21621 6953
rect 23293 6953 23305 6956
rect 23339 6953 23351 6987
rect 23293 6947 23351 6953
rect 23385 6987 23443 6993
rect 23385 6953 23397 6987
rect 23431 6984 23443 6987
rect 23658 6984 23664 6996
rect 23431 6956 23664 6984
rect 23431 6953 23443 6956
rect 23385 6947 23443 6953
rect 23658 6944 23664 6956
rect 23716 6944 23722 6996
rect 25038 6944 25044 6996
rect 25096 6984 25102 6996
rect 25317 6987 25375 6993
rect 25317 6984 25329 6987
rect 25096 6956 25329 6984
rect 25096 6944 25102 6956
rect 25317 6953 25329 6956
rect 25363 6984 25375 6987
rect 25590 6984 25596 6996
rect 25363 6956 25596 6984
rect 25363 6953 25375 6956
rect 25317 6947 25375 6953
rect 25590 6944 25596 6956
rect 25648 6944 25654 6996
rect 23566 6876 23572 6928
rect 23624 6916 23630 6928
rect 23624 6888 25728 6916
rect 23624 6876 23630 6888
rect 21821 6851 21879 6857
rect 21821 6817 21833 6851
rect 21867 6848 21879 6851
rect 23198 6848 23204 6860
rect 21867 6820 23204 6848
rect 21867 6817 21879 6820
rect 21821 6811 21879 6817
rect 23198 6808 23204 6820
rect 23256 6808 23262 6860
rect 23400 6820 23796 6848
rect 16393 6783 16451 6789
rect 16393 6749 16405 6783
rect 16439 6749 16451 6783
rect 16393 6743 16451 6749
rect 16408 6712 16436 6743
rect 18230 6740 18236 6792
rect 18288 6780 18294 6792
rect 18509 6783 18567 6789
rect 18509 6780 18521 6783
rect 18288 6752 18521 6780
rect 18288 6740 18294 6752
rect 18509 6749 18521 6752
rect 18555 6749 18567 6783
rect 18509 6743 18567 6749
rect 18690 6740 18696 6792
rect 18748 6780 18754 6792
rect 18969 6783 19027 6789
rect 18969 6780 18981 6783
rect 18748 6752 18981 6780
rect 18748 6740 18754 6752
rect 18969 6749 18981 6752
rect 19015 6749 19027 6783
rect 18969 6743 19027 6749
rect 21913 6783 21971 6789
rect 21913 6749 21925 6783
rect 21959 6780 21971 6783
rect 22186 6780 22192 6792
rect 21959 6752 22192 6780
rect 21959 6749 21971 6752
rect 21913 6743 21971 6749
rect 21818 6712 21824 6724
rect 16408 6684 16620 6712
rect 17894 6684 18276 6712
rect 21114 6684 21824 6712
rect 16592 6656 16620 6684
rect 18248 6656 18276 6684
rect 21818 6672 21824 6684
rect 21876 6672 21882 6724
rect 16574 6604 16580 6656
rect 16632 6604 16638 6656
rect 18230 6604 18236 6656
rect 18288 6604 18294 6656
rect 18782 6604 18788 6656
rect 18840 6604 18846 6656
rect 20073 6647 20131 6653
rect 20073 6613 20085 6647
rect 20119 6644 20131 6647
rect 21928 6644 21956 6743
rect 22186 6740 22192 6752
rect 22244 6740 22250 6792
rect 22557 6783 22615 6789
rect 22557 6749 22569 6783
rect 22603 6780 22615 6783
rect 23017 6783 23075 6789
rect 23017 6780 23029 6783
rect 22603 6752 23029 6780
rect 22603 6749 22615 6752
rect 22557 6743 22615 6749
rect 23017 6749 23029 6752
rect 23063 6749 23075 6783
rect 23017 6743 23075 6749
rect 23109 6783 23167 6789
rect 23109 6749 23121 6783
rect 23155 6780 23167 6783
rect 23400 6780 23428 6820
rect 23768 6792 23796 6820
rect 24946 6808 24952 6860
rect 25004 6808 25010 6860
rect 25700 6792 25728 6888
rect 23155 6752 23428 6780
rect 23155 6749 23167 6752
rect 23109 6743 23167 6749
rect 23474 6740 23480 6792
rect 23532 6780 23538 6792
rect 23569 6783 23627 6789
rect 23569 6780 23581 6783
rect 23532 6752 23581 6780
rect 23532 6740 23538 6752
rect 23569 6749 23581 6752
rect 23615 6749 23627 6783
rect 23569 6743 23627 6749
rect 23750 6740 23756 6792
rect 23808 6740 23814 6792
rect 23937 6783 23995 6789
rect 23937 6749 23949 6783
rect 23983 6780 23995 6783
rect 24397 6783 24455 6789
rect 24397 6780 24409 6783
rect 23983 6752 24409 6780
rect 23983 6749 23995 6752
rect 23937 6743 23995 6749
rect 24397 6749 24409 6752
rect 24443 6749 24455 6783
rect 24397 6743 24455 6749
rect 25409 6783 25467 6789
rect 25409 6749 25421 6783
rect 25455 6780 25467 6783
rect 25455 6752 25544 6780
rect 25455 6749 25467 6752
rect 25409 6743 25467 6749
rect 22370 6672 22376 6724
rect 22428 6712 22434 6724
rect 23661 6715 23719 6721
rect 23661 6712 23673 6715
rect 22428 6684 23673 6712
rect 22428 6672 22434 6684
rect 23661 6681 23673 6684
rect 23707 6681 23719 6715
rect 23661 6675 23719 6681
rect 25516 6656 25544 6752
rect 25682 6740 25688 6792
rect 25740 6740 25746 6792
rect 20119 6616 21956 6644
rect 20119 6613 20131 6616
rect 20073 6607 20131 6613
rect 22646 6604 22652 6656
rect 22704 6604 22710 6656
rect 23290 6604 23296 6656
rect 23348 6644 23354 6656
rect 25038 6644 25044 6656
rect 23348 6616 25044 6644
rect 23348 6604 23354 6616
rect 25038 6604 25044 6616
rect 25096 6604 25102 6656
rect 25130 6604 25136 6656
rect 25188 6604 25194 6656
rect 25498 6604 25504 6656
rect 25556 6604 25562 6656
rect 1104 6554 28888 6576
rect 1104 6502 5083 6554
rect 5135 6502 5147 6554
rect 5199 6502 5211 6554
rect 5263 6502 5275 6554
rect 5327 6502 5339 6554
rect 5391 6502 12029 6554
rect 12081 6502 12093 6554
rect 12145 6502 12157 6554
rect 12209 6502 12221 6554
rect 12273 6502 12285 6554
rect 12337 6502 18975 6554
rect 19027 6502 19039 6554
rect 19091 6502 19103 6554
rect 19155 6502 19167 6554
rect 19219 6502 19231 6554
rect 19283 6502 25921 6554
rect 25973 6502 25985 6554
rect 26037 6502 26049 6554
rect 26101 6502 26113 6554
rect 26165 6502 26177 6554
rect 26229 6502 28888 6554
rect 1104 6480 28888 6502
rect 20349 6443 20407 6449
rect 20349 6440 20361 6443
rect 18524 6412 19656 6440
rect 18230 6372 18236 6384
rect 18170 6344 18236 6372
rect 18230 6332 18236 6344
rect 18288 6372 18294 6384
rect 18524 6372 18552 6412
rect 19628 6372 19656 6412
rect 19996 6412 20361 6440
rect 19702 6372 19708 6384
rect 18288 6344 18552 6372
rect 19550 6344 19708 6372
rect 18288 6332 18294 6344
rect 19702 6332 19708 6344
rect 19760 6332 19766 6384
rect 19996 6381 20024 6412
rect 20349 6409 20361 6412
rect 20395 6409 20407 6443
rect 20349 6403 20407 6409
rect 22186 6400 22192 6452
rect 22244 6400 22250 6452
rect 22646 6400 22652 6452
rect 22704 6400 22710 6452
rect 23198 6400 23204 6452
rect 23256 6440 23262 6452
rect 23566 6440 23572 6452
rect 23256 6412 23572 6440
rect 23256 6400 23262 6412
rect 23566 6400 23572 6412
rect 23624 6400 23630 6452
rect 23750 6400 23756 6452
rect 23808 6440 23814 6452
rect 23845 6443 23903 6449
rect 23845 6440 23857 6443
rect 23808 6412 23857 6440
rect 23808 6400 23814 6412
rect 23845 6409 23857 6412
rect 23891 6409 23903 6443
rect 23845 6403 23903 6409
rect 19981 6375 20039 6381
rect 19981 6341 19993 6375
rect 20027 6341 20039 6375
rect 22204 6372 22232 6400
rect 22830 6372 22836 6384
rect 22204 6344 22836 6372
rect 19981 6335 20039 6341
rect 20530 6264 20536 6316
rect 20588 6264 20594 6316
rect 20714 6264 20720 6316
rect 20772 6304 20778 6316
rect 20993 6307 21051 6313
rect 20993 6304 21005 6307
rect 20772 6276 21005 6304
rect 20772 6264 20778 6276
rect 20993 6273 21005 6276
rect 21039 6273 21051 6307
rect 20993 6267 21051 6273
rect 21174 6264 21180 6316
rect 21232 6264 21238 6316
rect 22186 6264 22192 6316
rect 22244 6304 22250 6316
rect 22388 6313 22416 6344
rect 22830 6332 22836 6344
rect 22888 6332 22894 6384
rect 23109 6375 23167 6381
rect 23109 6341 23121 6375
rect 23155 6372 23167 6375
rect 24762 6372 24768 6384
rect 23155 6344 23888 6372
rect 23155 6341 23167 6344
rect 23109 6335 23167 6341
rect 23860 6316 23888 6344
rect 24044 6344 24768 6372
rect 24044 6316 24072 6344
rect 24762 6332 24768 6344
rect 24820 6332 24826 6384
rect 24946 6332 24952 6384
rect 25004 6332 25010 6384
rect 22281 6307 22339 6313
rect 22281 6304 22293 6307
rect 22244 6276 22293 6304
rect 22244 6264 22250 6276
rect 22281 6273 22293 6276
rect 22327 6273 22339 6307
rect 22281 6267 22339 6273
rect 22373 6307 22431 6313
rect 22373 6273 22385 6307
rect 22419 6273 22431 6307
rect 22373 6267 22431 6273
rect 23014 6264 23020 6316
rect 23072 6264 23078 6316
rect 23290 6264 23296 6316
rect 23348 6304 23354 6316
rect 23569 6307 23627 6313
rect 23569 6304 23581 6307
rect 23348 6276 23581 6304
rect 23348 6264 23354 6276
rect 23569 6273 23581 6276
rect 23615 6273 23627 6307
rect 23569 6267 23627 6273
rect 23753 6307 23811 6313
rect 23753 6273 23765 6307
rect 23799 6273 23811 6307
rect 23753 6267 23811 6273
rect 16574 6196 16580 6248
rect 16632 6236 16638 6248
rect 16669 6239 16727 6245
rect 16669 6236 16681 6239
rect 16632 6208 16681 6236
rect 16632 6196 16638 6208
rect 16669 6205 16681 6208
rect 16715 6205 16727 6239
rect 16669 6199 16727 6205
rect 16945 6239 17003 6245
rect 16945 6205 16957 6239
rect 16991 6236 17003 6239
rect 17402 6236 17408 6248
rect 16991 6208 17408 6236
rect 16991 6205 17003 6208
rect 16945 6199 17003 6205
rect 17402 6196 17408 6208
rect 17460 6196 17466 6248
rect 18417 6239 18475 6245
rect 18417 6205 18429 6239
rect 18463 6236 18475 6239
rect 19334 6236 19340 6248
rect 18463 6208 19340 6236
rect 18463 6205 18475 6208
rect 18417 6199 18475 6205
rect 19334 6196 19340 6208
rect 19392 6196 19398 6248
rect 20257 6239 20315 6245
rect 20257 6236 20269 6239
rect 20180 6208 20269 6236
rect 20180 6112 20208 6208
rect 20257 6205 20269 6208
rect 20303 6205 20315 6239
rect 23308 6236 23336 6264
rect 20257 6199 20315 6205
rect 22572 6208 23336 6236
rect 23385 6239 23443 6245
rect 21177 6171 21235 6177
rect 21177 6137 21189 6171
rect 21223 6168 21235 6171
rect 22370 6168 22376 6180
rect 21223 6140 22376 6168
rect 21223 6137 21235 6140
rect 21177 6131 21235 6137
rect 22370 6128 22376 6140
rect 22428 6128 22434 6180
rect 22572 6112 22600 6208
rect 23385 6205 23397 6239
rect 23431 6236 23443 6239
rect 23474 6236 23480 6248
rect 23431 6208 23480 6236
rect 23431 6205 23443 6208
rect 23385 6199 23443 6205
rect 23474 6196 23480 6208
rect 23532 6236 23538 6248
rect 23768 6236 23796 6267
rect 23842 6264 23848 6316
rect 23900 6264 23906 6316
rect 24026 6264 24032 6316
rect 24084 6264 24090 6316
rect 28258 6264 28264 6316
rect 28316 6264 28322 6316
rect 23532 6208 23796 6236
rect 23532 6196 23538 6208
rect 24210 6196 24216 6248
rect 24268 6196 24274 6248
rect 24486 6196 24492 6248
rect 24544 6196 24550 6248
rect 24578 6196 24584 6248
rect 24636 6236 24642 6248
rect 25498 6236 25504 6248
rect 24636 6208 25504 6236
rect 24636 6196 24642 6208
rect 25498 6196 25504 6208
rect 25556 6236 25562 6248
rect 25961 6239 26019 6245
rect 25961 6236 25973 6239
rect 25556 6208 25973 6236
rect 25556 6196 25562 6208
rect 25961 6205 25973 6208
rect 26007 6236 26019 6239
rect 26697 6239 26755 6245
rect 26697 6236 26709 6239
rect 26007 6208 26709 6236
rect 26007 6205 26019 6208
rect 25961 6199 26019 6205
rect 26697 6205 26709 6208
rect 26743 6205 26755 6239
rect 26697 6199 26755 6205
rect 28534 6196 28540 6248
rect 28592 6196 28598 6248
rect 26145 6171 26203 6177
rect 26145 6168 26157 6171
rect 25516 6140 26157 6168
rect 18509 6103 18567 6109
rect 18509 6069 18521 6103
rect 18555 6100 18567 6103
rect 19794 6100 19800 6112
rect 18555 6072 19800 6100
rect 18555 6069 18567 6072
rect 18509 6063 18567 6069
rect 19794 6060 19800 6072
rect 19852 6060 19858 6112
rect 20162 6060 20168 6112
rect 20220 6060 20226 6112
rect 22465 6103 22523 6109
rect 22465 6069 22477 6103
rect 22511 6100 22523 6103
rect 22554 6100 22560 6112
rect 22511 6072 22560 6100
rect 22511 6069 22523 6072
rect 22465 6063 22523 6069
rect 22554 6060 22560 6072
rect 22612 6060 22618 6112
rect 25038 6060 25044 6112
rect 25096 6100 25102 6112
rect 25516 6100 25544 6140
rect 26145 6137 26157 6140
rect 26191 6137 26203 6171
rect 26145 6131 26203 6137
rect 25096 6072 25544 6100
rect 25096 6060 25102 6072
rect 1104 6010 28888 6032
rect 1104 5958 4423 6010
rect 4475 5958 4487 6010
rect 4539 5958 4551 6010
rect 4603 5958 4615 6010
rect 4667 5958 4679 6010
rect 4731 5958 11369 6010
rect 11421 5958 11433 6010
rect 11485 5958 11497 6010
rect 11549 5958 11561 6010
rect 11613 5958 11625 6010
rect 11677 5958 18315 6010
rect 18367 5958 18379 6010
rect 18431 5958 18443 6010
rect 18495 5958 18507 6010
rect 18559 5958 18571 6010
rect 18623 5958 25261 6010
rect 25313 5958 25325 6010
rect 25377 5958 25389 6010
rect 25441 5958 25453 6010
rect 25505 5958 25517 6010
rect 25569 5958 28888 6010
rect 1104 5936 28888 5958
rect 19061 5899 19119 5905
rect 19061 5865 19073 5899
rect 19107 5896 19119 5899
rect 20530 5896 20536 5908
rect 19107 5868 20536 5896
rect 19107 5865 19119 5868
rect 19061 5859 19119 5865
rect 20530 5856 20536 5868
rect 20588 5856 20594 5908
rect 22738 5856 22744 5908
rect 22796 5896 22802 5908
rect 23477 5899 23535 5905
rect 23477 5896 23489 5899
rect 22796 5868 23489 5896
rect 22796 5856 22802 5868
rect 23477 5865 23489 5868
rect 23523 5865 23535 5899
rect 23477 5859 23535 5865
rect 24397 5899 24455 5905
rect 24397 5865 24409 5899
rect 24443 5896 24455 5899
rect 24486 5896 24492 5908
rect 24443 5868 24492 5896
rect 24443 5865 24455 5868
rect 24397 5859 24455 5865
rect 24486 5856 24492 5868
rect 24544 5856 24550 5908
rect 24578 5856 24584 5908
rect 24636 5856 24642 5908
rect 25038 5856 25044 5908
rect 25096 5856 25102 5908
rect 25130 5856 25136 5908
rect 25188 5856 25194 5908
rect 19334 5828 19340 5840
rect 17604 5800 19340 5828
rect 17604 5769 17632 5800
rect 19334 5788 19340 5800
rect 19392 5788 19398 5840
rect 17589 5763 17647 5769
rect 17589 5729 17601 5763
rect 17635 5729 17647 5763
rect 17589 5723 17647 5729
rect 18141 5763 18199 5769
rect 18141 5729 18153 5763
rect 18187 5760 18199 5763
rect 18601 5763 18659 5769
rect 18601 5760 18613 5763
rect 18187 5732 18613 5760
rect 18187 5729 18199 5732
rect 18141 5723 18199 5729
rect 18601 5729 18613 5732
rect 18647 5729 18659 5763
rect 18601 5723 18659 5729
rect 18693 5763 18751 5769
rect 18693 5729 18705 5763
rect 18739 5760 18751 5763
rect 19245 5763 19303 5769
rect 19245 5760 19257 5763
rect 18739 5732 19257 5760
rect 18739 5729 18751 5732
rect 18693 5723 18751 5729
rect 19245 5729 19257 5732
rect 19291 5729 19303 5763
rect 19245 5723 19303 5729
rect 19794 5720 19800 5772
rect 19852 5720 19858 5772
rect 20441 5763 20499 5769
rect 20441 5729 20453 5763
rect 20487 5760 20499 5763
rect 22005 5763 22063 5769
rect 22005 5760 22017 5763
rect 20487 5732 22017 5760
rect 20487 5729 20499 5732
rect 20441 5723 20499 5729
rect 22005 5729 22017 5732
rect 22051 5729 22063 5763
rect 23014 5760 23020 5772
rect 22005 5723 22063 5729
rect 22112 5732 23020 5760
rect 17862 5692 17868 5704
rect 17420 5664 17868 5692
rect 17420 5633 17448 5664
rect 17862 5652 17868 5664
rect 17920 5652 17926 5704
rect 18417 5695 18475 5701
rect 18417 5661 18429 5695
rect 18463 5692 18475 5695
rect 18877 5695 18935 5701
rect 18877 5692 18889 5695
rect 18463 5664 18889 5692
rect 18463 5661 18475 5664
rect 18417 5655 18475 5661
rect 18877 5661 18889 5664
rect 18923 5692 18935 5695
rect 20070 5692 20076 5704
rect 18923 5664 20076 5692
rect 18923 5661 18935 5664
rect 18877 5655 18935 5661
rect 20070 5652 20076 5664
rect 20128 5652 20134 5704
rect 20162 5652 20168 5704
rect 20220 5652 20226 5704
rect 21726 5692 21732 5704
rect 21574 5664 21732 5692
rect 21726 5652 21732 5664
rect 21784 5652 21790 5704
rect 17405 5627 17463 5633
rect 17405 5593 17417 5627
rect 17451 5593 17463 5627
rect 20180 5624 20208 5652
rect 22112 5636 22140 5732
rect 23014 5720 23020 5732
rect 23072 5760 23078 5772
rect 23293 5763 23351 5769
rect 23293 5760 23305 5763
rect 23072 5732 23305 5760
rect 23072 5720 23078 5732
rect 23293 5729 23305 5732
rect 23339 5760 23351 5763
rect 23934 5760 23940 5772
rect 23339 5732 23940 5760
rect 23339 5729 23351 5732
rect 23293 5723 23351 5729
rect 23934 5720 23940 5732
rect 23992 5720 23998 5772
rect 24596 5760 24624 5856
rect 25056 5828 25084 5856
rect 24688 5800 25084 5828
rect 24688 5769 24716 5800
rect 24504 5732 24624 5760
rect 24673 5763 24731 5769
rect 22190 5673 22248 5679
rect 22190 5639 22202 5673
rect 22236 5639 22248 5673
rect 22370 5652 22376 5704
rect 22428 5652 22434 5704
rect 22649 5695 22707 5701
rect 22649 5661 22661 5695
rect 22695 5692 22707 5695
rect 22741 5695 22799 5701
rect 22741 5692 22753 5695
rect 22695 5664 22753 5692
rect 22695 5661 22707 5664
rect 22649 5655 22707 5661
rect 22741 5661 22753 5664
rect 22787 5661 22799 5695
rect 22741 5655 22799 5661
rect 23658 5652 23664 5704
rect 23716 5652 23722 5704
rect 23750 5652 23756 5704
rect 23808 5652 23814 5704
rect 23842 5652 23848 5704
rect 23900 5692 23906 5704
rect 24504 5692 24532 5732
rect 24673 5729 24685 5763
rect 24719 5729 24731 5763
rect 24673 5723 24731 5729
rect 24762 5720 24768 5772
rect 24820 5720 24826 5772
rect 25041 5763 25099 5769
rect 25041 5729 25053 5763
rect 25087 5760 25099 5763
rect 25148 5760 25176 5856
rect 25682 5828 25688 5840
rect 25087 5732 25176 5760
rect 25424 5800 25688 5828
rect 25087 5729 25099 5732
rect 25041 5723 25099 5729
rect 23900 5664 24532 5692
rect 24581 5695 24639 5701
rect 23900 5652 23906 5664
rect 24581 5661 24593 5695
rect 24627 5661 24639 5695
rect 24780 5692 24808 5720
rect 25424 5701 25452 5800
rect 25682 5788 25688 5800
rect 25740 5788 25746 5840
rect 25133 5695 25191 5701
rect 25133 5692 25145 5695
rect 24780 5664 25145 5692
rect 24581 5655 24639 5661
rect 25133 5661 25145 5664
rect 25179 5661 25191 5695
rect 25133 5655 25191 5661
rect 25409 5695 25467 5701
rect 25409 5661 25421 5695
rect 25455 5661 25467 5695
rect 25409 5655 25467 5661
rect 22190 5636 22248 5639
rect 22094 5624 22100 5636
rect 17405 5587 17463 5593
rect 19812 5596 20208 5624
rect 21928 5596 22100 5624
rect 19812 5568 19840 5596
rect 16117 5559 16175 5565
rect 16117 5525 16129 5559
rect 16163 5556 16175 5559
rect 16574 5556 16580 5568
rect 16163 5528 16580 5556
rect 16163 5525 16175 5528
rect 16117 5519 16175 5525
rect 16574 5516 16580 5528
rect 16632 5516 16638 5568
rect 17954 5516 17960 5568
rect 18012 5556 18018 5568
rect 18233 5559 18291 5565
rect 18233 5556 18245 5559
rect 18012 5528 18245 5556
rect 18012 5516 18018 5528
rect 18233 5525 18245 5528
rect 18279 5525 18291 5559
rect 18233 5519 18291 5525
rect 19794 5516 19800 5568
rect 19852 5516 19858 5568
rect 21928 5565 21956 5596
rect 22094 5584 22100 5596
rect 22152 5584 22158 5636
rect 22186 5584 22192 5636
rect 22244 5584 22250 5636
rect 22278 5584 22284 5636
rect 22336 5584 22342 5636
rect 22462 5584 22468 5636
rect 22520 5633 22526 5636
rect 22520 5627 22549 5633
rect 22537 5593 22549 5627
rect 22520 5587 22549 5593
rect 22520 5584 22526 5587
rect 24302 5584 24308 5636
rect 24360 5624 24366 5636
rect 24596 5624 24624 5655
rect 25590 5652 25596 5704
rect 25648 5652 25654 5704
rect 24360 5596 25176 5624
rect 24360 5584 24366 5596
rect 21913 5559 21971 5565
rect 21913 5525 21925 5559
rect 21959 5525 21971 5559
rect 25148 5556 25176 5596
rect 25317 5559 25375 5565
rect 25317 5556 25329 5559
rect 25148 5528 25329 5556
rect 21913 5519 21971 5525
rect 25317 5525 25329 5528
rect 25363 5525 25375 5559
rect 25317 5519 25375 5525
rect 1104 5466 28888 5488
rect 1104 5414 5083 5466
rect 5135 5414 5147 5466
rect 5199 5414 5211 5466
rect 5263 5414 5275 5466
rect 5327 5414 5339 5466
rect 5391 5414 12029 5466
rect 12081 5414 12093 5466
rect 12145 5414 12157 5466
rect 12209 5414 12221 5466
rect 12273 5414 12285 5466
rect 12337 5414 18975 5466
rect 19027 5414 19039 5466
rect 19091 5414 19103 5466
rect 19155 5414 19167 5466
rect 19219 5414 19231 5466
rect 19283 5414 25921 5466
rect 25973 5414 25985 5466
rect 26037 5414 26049 5466
rect 26101 5414 26113 5466
rect 26165 5414 26177 5466
rect 26229 5414 28888 5466
rect 1104 5392 28888 5414
rect 19705 5355 19763 5361
rect 16960 5324 18828 5352
rect 16960 5293 16988 5324
rect 18800 5296 18828 5324
rect 19705 5321 19717 5355
rect 19751 5352 19763 5355
rect 20257 5355 20315 5361
rect 19751 5324 19840 5352
rect 19751 5321 19763 5324
rect 19705 5315 19763 5321
rect 16945 5287 17003 5293
rect 16945 5253 16957 5287
rect 16991 5253 17003 5287
rect 16945 5247 17003 5253
rect 18782 5244 18788 5296
rect 18840 5244 18846 5296
rect 19812 5293 19840 5324
rect 20257 5321 20269 5355
rect 20303 5352 20315 5355
rect 21910 5352 21916 5364
rect 20303 5324 21916 5352
rect 20303 5321 20315 5324
rect 20257 5315 20315 5321
rect 21910 5312 21916 5324
rect 21968 5312 21974 5364
rect 22094 5312 22100 5364
rect 22152 5312 22158 5364
rect 22186 5312 22192 5364
rect 22244 5352 22250 5364
rect 22465 5355 22523 5361
rect 22465 5352 22477 5355
rect 22244 5324 22477 5352
rect 22244 5312 22250 5324
rect 22465 5321 22477 5324
rect 22511 5321 22523 5355
rect 22465 5315 22523 5321
rect 22922 5312 22928 5364
rect 22980 5352 22986 5364
rect 23198 5352 23204 5364
rect 22980 5324 23204 5352
rect 22980 5312 22986 5324
rect 23198 5312 23204 5324
rect 23256 5312 23262 5364
rect 23385 5355 23443 5361
rect 23385 5321 23397 5355
rect 23431 5321 23443 5355
rect 23750 5352 23756 5364
rect 23385 5315 23443 5321
rect 23676 5324 23756 5352
rect 19797 5287 19855 5293
rect 19797 5253 19809 5287
rect 19843 5253 19855 5287
rect 19797 5247 19855 5253
rect 20548 5256 22048 5284
rect 16574 5108 16580 5160
rect 16632 5148 16638 5160
rect 16669 5151 16727 5157
rect 16669 5148 16681 5151
rect 16632 5120 16681 5148
rect 16632 5108 16638 5120
rect 16669 5117 16681 5120
rect 16715 5117 16727 5151
rect 18064 5148 18092 5202
rect 18230 5176 18236 5228
rect 18288 5216 18294 5228
rect 19245 5219 19303 5225
rect 19245 5216 19257 5219
rect 18288 5188 19257 5216
rect 18288 5176 18294 5188
rect 19245 5185 19257 5188
rect 19291 5185 19303 5219
rect 19245 5179 19303 5185
rect 19426 5176 19432 5228
rect 19484 5216 19490 5228
rect 19521 5219 19579 5225
rect 19521 5216 19533 5219
rect 19484 5188 19533 5216
rect 19484 5176 19490 5188
rect 19521 5185 19533 5188
rect 19567 5185 19579 5219
rect 19521 5179 19579 5185
rect 19886 5176 19892 5228
rect 19944 5216 19950 5228
rect 20073 5219 20131 5225
rect 20073 5216 20085 5219
rect 19944 5188 20085 5216
rect 19944 5176 19950 5188
rect 20073 5185 20085 5188
rect 20119 5185 20131 5219
rect 20073 5179 20131 5185
rect 20254 5176 20260 5228
rect 20312 5216 20318 5228
rect 20548 5225 20576 5256
rect 20533 5219 20591 5225
rect 20533 5216 20545 5219
rect 20312 5188 20545 5216
rect 20312 5176 20318 5188
rect 20533 5185 20545 5188
rect 20579 5185 20591 5219
rect 20990 5216 20996 5228
rect 20533 5179 20591 5185
rect 20640 5188 20996 5216
rect 18322 5148 18328 5160
rect 18064 5120 18328 5148
rect 16669 5111 16727 5117
rect 18322 5108 18328 5120
rect 18380 5108 18386 5160
rect 18417 5151 18475 5157
rect 18417 5117 18429 5151
rect 18463 5148 18475 5151
rect 19061 5151 19119 5157
rect 19061 5148 19073 5151
rect 18463 5120 19073 5148
rect 18463 5117 18475 5120
rect 18417 5111 18475 5117
rect 19061 5117 19073 5120
rect 19107 5148 19119 5151
rect 19337 5151 19395 5157
rect 19337 5148 19349 5151
rect 19107 5120 19349 5148
rect 19107 5117 19119 5120
rect 19061 5111 19119 5117
rect 19337 5117 19349 5120
rect 19383 5117 19395 5151
rect 19337 5111 19395 5117
rect 19981 5151 20039 5157
rect 19981 5117 19993 5151
rect 20027 5148 20039 5151
rect 20640 5148 20668 5188
rect 20990 5176 20996 5188
rect 21048 5216 21054 5228
rect 21361 5219 21419 5225
rect 21361 5216 21373 5219
rect 21048 5188 21373 5216
rect 21048 5176 21054 5188
rect 21361 5185 21373 5188
rect 21407 5185 21419 5219
rect 21361 5179 21419 5185
rect 21634 5176 21640 5228
rect 21692 5216 21698 5228
rect 21821 5219 21879 5225
rect 21821 5216 21833 5219
rect 21692 5188 21833 5216
rect 21692 5176 21698 5188
rect 21821 5185 21833 5188
rect 21867 5185 21879 5219
rect 21821 5179 21879 5185
rect 20027 5120 20668 5148
rect 20717 5151 20775 5157
rect 20027 5117 20039 5120
rect 19981 5111 20039 5117
rect 20717 5117 20729 5151
rect 20763 5148 20775 5151
rect 20809 5151 20867 5157
rect 20809 5148 20821 5151
rect 20763 5120 20821 5148
rect 20763 5117 20775 5120
rect 20717 5111 20775 5117
rect 20809 5117 20821 5120
rect 20855 5117 20867 5151
rect 20809 5111 20867 5117
rect 18340 5080 18368 5108
rect 18966 5080 18972 5092
rect 18340 5052 18972 5080
rect 18966 5040 18972 5052
rect 19024 5040 19030 5092
rect 18046 4972 18052 5024
rect 18104 5012 18110 5024
rect 18509 5015 18567 5021
rect 18509 5012 18521 5015
rect 18104 4984 18521 5012
rect 18104 4972 18110 4984
rect 18509 4981 18521 4984
rect 18555 4981 18567 5015
rect 18509 4975 18567 4981
rect 19334 4972 19340 5024
rect 19392 4972 19398 5024
rect 19702 4972 19708 5024
rect 19760 5012 19766 5024
rect 19797 5015 19855 5021
rect 19797 5012 19809 5015
rect 19760 4984 19809 5012
rect 19760 4972 19766 4984
rect 19797 4981 19809 4984
rect 19843 4981 19855 5015
rect 19797 4975 19855 4981
rect 20346 4972 20352 5024
rect 20404 4972 20410 5024
rect 21836 5012 21864 5179
rect 22020 5089 22048 5256
rect 22112 5216 22140 5312
rect 22278 5244 22284 5296
rect 22336 5284 22342 5296
rect 23400 5284 23428 5315
rect 22336 5256 23428 5284
rect 22336 5244 22342 5256
rect 22465 5219 22523 5225
rect 22465 5216 22477 5219
rect 22112 5188 22477 5216
rect 22465 5185 22477 5188
rect 22511 5185 22523 5219
rect 22465 5179 22523 5185
rect 22557 5219 22615 5225
rect 22557 5185 22569 5219
rect 22603 5185 22615 5219
rect 22557 5179 22615 5185
rect 22741 5219 22799 5225
rect 22741 5185 22753 5219
rect 22787 5216 22799 5219
rect 22922 5216 22928 5228
rect 22787 5188 22928 5216
rect 22787 5185 22799 5188
rect 22741 5179 22799 5185
rect 22005 5083 22063 5089
rect 22005 5049 22017 5083
rect 22051 5080 22063 5083
rect 22462 5080 22468 5092
rect 22051 5052 22468 5080
rect 22051 5049 22063 5052
rect 22005 5043 22063 5049
rect 22462 5040 22468 5052
rect 22520 5040 22526 5092
rect 22278 5012 22284 5024
rect 21836 4984 22284 5012
rect 22278 4972 22284 4984
rect 22336 4972 22342 5024
rect 22572 5012 22600 5179
rect 22922 5176 22928 5188
rect 22980 5176 22986 5228
rect 23676 5225 23704 5324
rect 23750 5312 23756 5324
rect 23808 5352 23814 5364
rect 23808 5324 25912 5352
rect 23808 5312 23814 5324
rect 25225 5287 25283 5293
rect 25225 5284 25237 5287
rect 24136 5256 25237 5284
rect 23109 5219 23167 5225
rect 23109 5216 23121 5219
rect 23032 5188 23121 5216
rect 23032 5092 23060 5188
rect 23109 5185 23121 5188
rect 23155 5216 23167 5219
rect 23569 5219 23627 5225
rect 23569 5216 23581 5219
rect 23155 5188 23581 5216
rect 23155 5185 23167 5188
rect 23109 5179 23167 5185
rect 23569 5185 23581 5188
rect 23615 5185 23627 5219
rect 23569 5179 23627 5185
rect 23661 5219 23719 5225
rect 23661 5185 23673 5219
rect 23707 5185 23719 5219
rect 23661 5179 23719 5185
rect 23293 5151 23351 5157
rect 23293 5117 23305 5151
rect 23339 5148 23351 5151
rect 23676 5148 23704 5179
rect 23750 5176 23756 5228
rect 23808 5176 23814 5228
rect 23845 5219 23903 5225
rect 23845 5185 23857 5219
rect 23891 5216 23903 5219
rect 23934 5216 23940 5228
rect 23891 5188 23940 5216
rect 23891 5185 23903 5188
rect 23845 5179 23903 5185
rect 23934 5176 23940 5188
rect 23992 5176 23998 5228
rect 24136 5225 24164 5256
rect 25225 5253 25237 5256
rect 25271 5253 25283 5287
rect 25225 5247 25283 5253
rect 24121 5219 24179 5225
rect 24121 5185 24133 5219
rect 24167 5185 24179 5219
rect 24121 5179 24179 5185
rect 24302 5176 24308 5228
rect 24360 5176 24366 5228
rect 24397 5219 24455 5225
rect 24397 5185 24409 5219
rect 24443 5185 24455 5219
rect 24397 5179 24455 5185
rect 24489 5219 24547 5225
rect 24489 5185 24501 5219
rect 24535 5216 24547 5219
rect 24765 5219 24823 5225
rect 24535 5188 24624 5216
rect 24535 5185 24547 5188
rect 24489 5179 24547 5185
rect 24412 5148 24440 5179
rect 23339 5120 23704 5148
rect 24320 5120 24440 5148
rect 23339 5117 23351 5120
rect 23293 5111 23351 5117
rect 23014 5040 23020 5092
rect 23072 5080 23078 5092
rect 24320 5080 24348 5120
rect 23072 5052 24348 5080
rect 24596 5080 24624 5188
rect 24765 5185 24777 5219
rect 24811 5185 24823 5219
rect 24765 5179 24823 5185
rect 24780 5148 24808 5179
rect 24854 5176 24860 5228
rect 24912 5216 24918 5228
rect 24949 5219 25007 5225
rect 24949 5216 24961 5219
rect 24912 5188 24961 5216
rect 24912 5176 24918 5188
rect 24949 5185 24961 5188
rect 24995 5216 25007 5219
rect 25590 5216 25596 5228
rect 24995 5188 25596 5216
rect 24995 5185 25007 5188
rect 24949 5179 25007 5185
rect 25590 5176 25596 5188
rect 25648 5176 25654 5228
rect 25682 5176 25688 5228
rect 25740 5176 25746 5228
rect 25700 5148 25728 5176
rect 25884 5157 25912 5324
rect 24780 5120 25728 5148
rect 25869 5151 25927 5157
rect 25869 5117 25881 5151
rect 25915 5148 25927 5151
rect 25915 5120 26188 5148
rect 25915 5117 25927 5120
rect 25869 5111 25927 5117
rect 24765 5083 24823 5089
rect 24765 5080 24777 5083
rect 24596 5052 24777 5080
rect 23072 5040 23078 5052
rect 24765 5049 24777 5052
rect 24811 5049 24823 5083
rect 24765 5043 24823 5049
rect 26160 5024 26188 5120
rect 23750 5012 23756 5024
rect 22572 4984 23756 5012
rect 23750 4972 23756 4984
rect 23808 4972 23814 5024
rect 24670 4972 24676 5024
rect 24728 4972 24734 5024
rect 26142 4972 26148 5024
rect 26200 4972 26206 5024
rect 1104 4922 28888 4944
rect 1104 4870 4423 4922
rect 4475 4870 4487 4922
rect 4539 4870 4551 4922
rect 4603 4870 4615 4922
rect 4667 4870 4679 4922
rect 4731 4870 11369 4922
rect 11421 4870 11433 4922
rect 11485 4870 11497 4922
rect 11549 4870 11561 4922
rect 11613 4870 11625 4922
rect 11677 4870 18315 4922
rect 18367 4870 18379 4922
rect 18431 4870 18443 4922
rect 18495 4870 18507 4922
rect 18559 4870 18571 4922
rect 18623 4870 25261 4922
rect 25313 4870 25325 4922
rect 25377 4870 25389 4922
rect 25441 4870 25453 4922
rect 25505 4870 25517 4922
rect 25569 4870 28888 4922
rect 1104 4848 28888 4870
rect 17402 4768 17408 4820
rect 17460 4808 17466 4820
rect 17773 4811 17831 4817
rect 17773 4808 17785 4811
rect 17460 4780 17785 4808
rect 17460 4768 17466 4780
rect 17773 4777 17785 4780
rect 17819 4777 17831 4811
rect 17773 4771 17831 4777
rect 18230 4768 18236 4820
rect 18288 4768 18294 4820
rect 18693 4811 18751 4817
rect 18693 4777 18705 4811
rect 18739 4808 18751 4811
rect 19334 4808 19340 4820
rect 18739 4780 19340 4808
rect 18739 4777 18751 4780
rect 18693 4771 18751 4777
rect 19334 4768 19340 4780
rect 19392 4768 19398 4820
rect 20990 4768 20996 4820
rect 21048 4768 21054 4820
rect 22278 4768 22284 4820
rect 22336 4808 22342 4820
rect 23290 4808 23296 4820
rect 22336 4780 23296 4808
rect 22336 4768 22342 4780
rect 23290 4768 23296 4780
rect 23348 4808 23354 4820
rect 24026 4808 24032 4820
rect 23348 4780 24032 4808
rect 23348 4768 23354 4780
rect 24026 4768 24032 4780
rect 24084 4768 24090 4820
rect 26142 4768 26148 4820
rect 26200 4768 26206 4820
rect 15841 4675 15899 4681
rect 15841 4641 15853 4675
rect 15887 4672 15899 4675
rect 16574 4672 16580 4684
rect 15887 4644 16580 4672
rect 15887 4641 15899 4644
rect 15841 4635 15899 4641
rect 16574 4632 16580 4644
rect 16632 4632 16638 4684
rect 17589 4675 17647 4681
rect 17589 4641 17601 4675
rect 17635 4672 17647 4675
rect 18141 4675 18199 4681
rect 18141 4672 18153 4675
rect 17635 4644 18153 4672
rect 17635 4641 17647 4644
rect 17589 4635 17647 4641
rect 18141 4641 18153 4644
rect 18187 4672 18199 4675
rect 18248 4672 18276 4768
rect 18874 4700 18880 4752
rect 18932 4740 18938 4752
rect 18969 4743 19027 4749
rect 18969 4740 18981 4743
rect 18932 4712 18981 4740
rect 18932 4700 18938 4712
rect 18969 4709 18981 4712
rect 19015 4709 19027 4743
rect 18969 4703 19027 4709
rect 21468 4712 23060 4740
rect 18187 4644 18276 4672
rect 18984 4644 20668 4672
rect 18187 4641 18199 4644
rect 18141 4635 18199 4641
rect 18984 4616 19012 4644
rect 17954 4564 17960 4616
rect 18012 4564 18018 4616
rect 18782 4564 18788 4616
rect 18840 4564 18846 4616
rect 18966 4564 18972 4616
rect 19024 4564 19030 4616
rect 19245 4607 19303 4613
rect 19245 4573 19257 4607
rect 19291 4573 19303 4607
rect 20640 4590 20668 4644
rect 21468 4616 21496 4712
rect 21560 4644 22784 4672
rect 19245 4567 19303 4573
rect 16114 4496 16120 4548
rect 16172 4496 16178 4548
rect 18984 4536 19012 4564
rect 17342 4508 19012 4536
rect 17972 4480 18000 4508
rect 17954 4428 17960 4480
rect 18012 4428 18018 4480
rect 19260 4468 19288 4567
rect 21266 4564 21272 4616
rect 21324 4564 21330 4616
rect 21450 4564 21456 4616
rect 21508 4564 21514 4616
rect 21560 4613 21588 4644
rect 22756 4616 22784 4644
rect 21545 4607 21603 4613
rect 21545 4573 21557 4607
rect 21591 4573 21603 4607
rect 21545 4567 21603 4573
rect 21729 4607 21787 4613
rect 21729 4573 21741 4607
rect 21775 4604 21787 4607
rect 22097 4607 22155 4613
rect 22097 4604 22109 4607
rect 21775 4576 22109 4604
rect 21775 4573 21787 4576
rect 21729 4567 21787 4573
rect 22097 4573 22109 4576
rect 22143 4604 22155 4607
rect 22143 4576 22197 4604
rect 22143 4573 22155 4576
rect 22097 4567 22155 4573
rect 19518 4496 19524 4548
rect 19576 4496 19582 4548
rect 19610 4496 19616 4548
rect 19668 4536 19674 4548
rect 19668 4508 19932 4536
rect 19668 4496 19674 4508
rect 19794 4468 19800 4480
rect 19260 4440 19800 4468
rect 19794 4428 19800 4440
rect 19852 4428 19858 4480
rect 19904 4468 19932 4508
rect 21085 4471 21143 4477
rect 21085 4468 21097 4471
rect 19904 4440 21097 4468
rect 21085 4437 21097 4440
rect 21131 4437 21143 4471
rect 21085 4431 21143 4437
rect 21542 4428 21548 4480
rect 21600 4468 21606 4480
rect 21744 4468 21772 4567
rect 22112 4536 22140 4567
rect 22738 4564 22744 4616
rect 22796 4564 22802 4616
rect 22830 4536 22836 4548
rect 22112 4508 22836 4536
rect 22830 4496 22836 4508
rect 22888 4496 22894 4548
rect 23032 4545 23060 4712
rect 24210 4632 24216 4684
rect 24268 4672 24274 4684
rect 24397 4675 24455 4681
rect 24397 4672 24409 4675
rect 24268 4644 24409 4672
rect 24268 4632 24274 4644
rect 24397 4641 24409 4644
rect 24443 4641 24455 4675
rect 24397 4635 24455 4641
rect 24670 4632 24676 4684
rect 24728 4632 24734 4684
rect 23661 4607 23719 4613
rect 23661 4573 23673 4607
rect 23707 4573 23719 4607
rect 23661 4567 23719 4573
rect 23017 4539 23075 4545
rect 23017 4505 23029 4539
rect 23063 4536 23075 4539
rect 23106 4536 23112 4548
rect 23063 4508 23112 4536
rect 23063 4505 23075 4508
rect 23017 4499 23075 4505
rect 23106 4496 23112 4508
rect 23164 4496 23170 4548
rect 23676 4536 23704 4567
rect 24946 4536 24952 4548
rect 23676 4508 24952 4536
rect 24946 4496 24952 4508
rect 25004 4496 25010 4548
rect 25130 4496 25136 4548
rect 25188 4496 25194 4548
rect 21600 4440 21772 4468
rect 21600 4428 21606 4440
rect 21910 4428 21916 4480
rect 21968 4428 21974 4480
rect 22646 4428 22652 4480
rect 22704 4428 22710 4480
rect 22922 4428 22928 4480
rect 22980 4468 22986 4480
rect 23290 4468 23296 4480
rect 22980 4440 23296 4468
rect 22980 4428 22986 4440
rect 23290 4428 23296 4440
rect 23348 4428 23354 4480
rect 23474 4428 23480 4480
rect 23532 4468 23538 4480
rect 23569 4471 23627 4477
rect 23569 4468 23581 4471
rect 23532 4440 23581 4468
rect 23532 4428 23538 4440
rect 23569 4437 23581 4440
rect 23615 4437 23627 4471
rect 23569 4431 23627 4437
rect 1104 4378 28888 4400
rect 1104 4326 5083 4378
rect 5135 4326 5147 4378
rect 5199 4326 5211 4378
rect 5263 4326 5275 4378
rect 5327 4326 5339 4378
rect 5391 4326 12029 4378
rect 12081 4326 12093 4378
rect 12145 4326 12157 4378
rect 12209 4326 12221 4378
rect 12273 4326 12285 4378
rect 12337 4326 18975 4378
rect 19027 4326 19039 4378
rect 19091 4326 19103 4378
rect 19155 4326 19167 4378
rect 19219 4326 19231 4378
rect 19283 4326 25921 4378
rect 25973 4326 25985 4378
rect 26037 4326 26049 4378
rect 26101 4326 26113 4378
rect 26165 4326 26177 4378
rect 26229 4326 28888 4378
rect 1104 4304 28888 4326
rect 16114 4224 16120 4276
rect 16172 4264 16178 4276
rect 16301 4267 16359 4273
rect 16301 4264 16313 4267
rect 16172 4236 16313 4264
rect 16172 4224 16178 4236
rect 16301 4233 16313 4236
rect 16347 4233 16359 4267
rect 16301 4227 16359 4233
rect 19429 4267 19487 4273
rect 19429 4233 19441 4267
rect 19475 4264 19487 4267
rect 19518 4264 19524 4276
rect 19475 4236 19524 4264
rect 19475 4233 19487 4236
rect 19429 4227 19487 4233
rect 19518 4224 19524 4236
rect 19576 4224 19582 4276
rect 20346 4224 20352 4276
rect 20404 4224 20410 4276
rect 21542 4224 21548 4276
rect 21600 4224 21606 4276
rect 21910 4224 21916 4276
rect 21968 4264 21974 4276
rect 21968 4236 22140 4264
rect 21968 4224 21974 4236
rect 20364 4196 20392 4224
rect 21726 4196 21732 4208
rect 17420 4168 17816 4196
rect 16485 4131 16543 4137
rect 16485 4097 16497 4131
rect 16531 4128 16543 4131
rect 17126 4128 17132 4140
rect 16531 4100 17132 4128
rect 16531 4097 16543 4100
rect 16485 4091 16543 4097
rect 17126 4088 17132 4100
rect 17184 4088 17190 4140
rect 17420 4137 17448 4168
rect 17405 4131 17463 4137
rect 17405 4097 17417 4131
rect 17451 4097 17463 4131
rect 17788 4126 17816 4168
rect 17972 4168 19564 4196
rect 17865 4132 17923 4137
rect 17972 4132 18000 4168
rect 17865 4131 18000 4132
rect 17865 4126 17877 4131
rect 17788 4098 17877 4126
rect 17405 4091 17463 4097
rect 17865 4097 17877 4098
rect 17911 4104 18000 4131
rect 17911 4097 17923 4104
rect 17865 4091 17923 4097
rect 18966 4088 18972 4140
rect 19024 4088 19030 4140
rect 19168 4137 19196 4168
rect 19153 4131 19211 4137
rect 19153 4097 19165 4131
rect 19199 4128 19211 4131
rect 19199 4100 19233 4128
rect 19199 4097 19211 4100
rect 19153 4091 19211 4097
rect 19334 4088 19340 4140
rect 19392 4088 19398 4140
rect 19426 4088 19432 4140
rect 19484 4088 19490 4140
rect 17589 4063 17647 4069
rect 17589 4029 17601 4063
rect 17635 4029 17647 4063
rect 17589 4023 17647 4029
rect 17681 4063 17739 4069
rect 17681 4029 17693 4063
rect 17727 4060 17739 4063
rect 18046 4060 18052 4072
rect 17727 4032 18052 4060
rect 17727 4029 17739 4032
rect 17681 4023 17739 4029
rect 17604 3992 17632 4023
rect 18046 4020 18052 4032
rect 18104 4020 18110 4072
rect 18690 4020 18696 4072
rect 18748 4020 18754 4072
rect 18877 4063 18935 4069
rect 18877 4029 18889 4063
rect 18923 4060 18935 4063
rect 19444 4060 19472 4088
rect 18923 4032 19472 4060
rect 18923 4029 18935 4032
rect 18877 4023 18935 4029
rect 18233 3995 18291 4001
rect 18233 3992 18245 3995
rect 17604 3964 18245 3992
rect 18233 3961 18245 3964
rect 18279 3961 18291 3995
rect 18233 3955 18291 3961
rect 17221 3927 17279 3933
rect 17221 3893 17233 3927
rect 17267 3924 17279 3927
rect 17402 3924 17408 3936
rect 17267 3896 17408 3924
rect 17267 3893 17279 3896
rect 17221 3887 17279 3893
rect 17402 3884 17408 3896
rect 17460 3884 17466 3936
rect 18049 3927 18107 3933
rect 18049 3893 18061 3927
rect 18095 3924 18107 3927
rect 18708 3924 18736 4020
rect 18095 3896 18736 3924
rect 19536 3924 19564 4168
rect 19628 4168 20392 4196
rect 21298 4168 21732 4196
rect 19628 4137 19656 4168
rect 21726 4156 21732 4168
rect 21784 4156 21790 4208
rect 22112 4205 22140 4236
rect 22462 4224 22468 4276
rect 22520 4224 22526 4276
rect 22557 4267 22615 4273
rect 22557 4233 22569 4267
rect 22603 4264 22615 4267
rect 23014 4264 23020 4276
rect 22603 4236 23020 4264
rect 22603 4233 22615 4236
rect 22557 4227 22615 4233
rect 23014 4224 23020 4236
rect 23072 4264 23078 4276
rect 23566 4264 23572 4276
rect 23072 4236 23572 4264
rect 23072 4224 23078 4236
rect 23566 4224 23572 4236
rect 23624 4224 23630 4276
rect 23937 4267 23995 4273
rect 23937 4233 23949 4267
rect 23983 4264 23995 4267
rect 24026 4264 24032 4276
rect 23983 4236 24032 4264
rect 23983 4233 23995 4236
rect 23937 4227 23995 4233
rect 24026 4224 24032 4236
rect 24084 4224 24090 4276
rect 24946 4224 24952 4276
rect 25004 4224 25010 4276
rect 22097 4199 22155 4205
rect 22097 4165 22109 4199
rect 22143 4165 22155 4199
rect 22097 4159 22155 4165
rect 22186 4156 22192 4208
rect 22244 4156 22250 4208
rect 22327 4199 22385 4205
rect 22327 4165 22339 4199
rect 22373 4196 22385 4199
rect 22480 4196 22508 4224
rect 22373 4168 22508 4196
rect 22741 4199 22799 4205
rect 22373 4165 22385 4168
rect 22327 4159 22385 4165
rect 22741 4165 22753 4199
rect 22787 4196 22799 4199
rect 22787 4168 23152 4196
rect 22787 4165 22799 4168
rect 22741 4159 22799 4165
rect 23124 4140 23152 4168
rect 23492 4168 23977 4196
rect 19613 4131 19671 4137
rect 19613 4097 19625 4131
rect 19659 4097 19671 4131
rect 19613 4091 19671 4097
rect 22005 4131 22063 4137
rect 22005 4097 22017 4131
rect 22051 4097 22063 4131
rect 22005 4091 22063 4097
rect 22465 4131 22523 4137
rect 22465 4097 22477 4131
rect 22511 4128 22523 4131
rect 22646 4128 22652 4140
rect 22511 4100 22652 4128
rect 22511 4097 22523 4100
rect 22465 4091 22523 4097
rect 19794 4020 19800 4072
rect 19852 4020 19858 4072
rect 20073 4063 20131 4069
rect 20073 4029 20085 4063
rect 20119 4060 20131 4063
rect 21821 4063 21879 4069
rect 21821 4060 21833 4063
rect 20119 4032 21833 4060
rect 20119 4029 20131 4032
rect 20073 4023 20131 4029
rect 21821 4029 21833 4032
rect 21867 4029 21879 4063
rect 22020 4060 22048 4091
rect 22646 4088 22652 4100
rect 22704 4088 22710 4140
rect 22830 4088 22836 4140
rect 22888 4088 22894 4140
rect 22925 4131 22983 4137
rect 22925 4097 22937 4131
rect 22971 4128 22983 4131
rect 23014 4128 23020 4140
rect 22971 4100 23020 4128
rect 22971 4097 22983 4100
rect 22925 4091 22983 4097
rect 23014 4088 23020 4100
rect 23072 4088 23078 4140
rect 23106 4088 23112 4140
rect 23164 4128 23170 4140
rect 23492 4137 23520 4168
rect 23201 4131 23259 4137
rect 23201 4128 23213 4131
rect 23164 4100 23213 4128
rect 23164 4088 23170 4100
rect 23201 4097 23213 4100
rect 23247 4097 23259 4131
rect 23201 4091 23259 4097
rect 23477 4131 23535 4137
rect 23477 4097 23489 4131
rect 23523 4097 23535 4131
rect 23477 4091 23535 4097
rect 22848 4060 22876 4088
rect 23293 4063 23351 4069
rect 23293 4060 23305 4063
rect 22020 4032 22094 4060
rect 22848 4032 23305 4060
rect 21821 4023 21879 4029
rect 22066 3992 22094 4032
rect 23293 4029 23305 4032
rect 23339 4029 23351 4063
rect 23293 4023 23351 4029
rect 22922 3992 22928 4004
rect 22066 3964 22928 3992
rect 22922 3952 22928 3964
rect 22980 3952 22986 4004
rect 23109 3995 23167 4001
rect 23109 3961 23121 3995
rect 23155 3992 23167 3995
rect 23492 3992 23520 4091
rect 23566 4088 23572 4140
rect 23624 4088 23630 4140
rect 23949 4137 23977 4168
rect 23934 4131 23992 4137
rect 23934 4097 23946 4131
rect 23980 4128 23992 4131
rect 23980 4100 25636 4128
rect 23980 4097 23992 4100
rect 23934 4091 23992 4097
rect 23584 4060 23612 4088
rect 24305 4063 24363 4069
rect 24305 4060 24317 4063
rect 23584 4032 24317 4060
rect 24305 4029 24317 4032
rect 24351 4029 24363 4063
rect 24305 4023 24363 4029
rect 24397 4063 24455 4069
rect 24397 4029 24409 4063
rect 24443 4060 24455 4063
rect 24762 4060 24768 4072
rect 24443 4032 24768 4060
rect 24443 4029 24455 4032
rect 24397 4023 24455 4029
rect 24762 4020 24768 4032
rect 24820 4020 24826 4072
rect 25608 4069 25636 4100
rect 25593 4063 25651 4069
rect 25593 4029 25605 4063
rect 25639 4060 25651 4063
rect 26142 4060 26148 4072
rect 25639 4032 26148 4060
rect 25639 4029 25651 4032
rect 25593 4023 25651 4029
rect 26142 4020 26148 4032
rect 26200 4020 26206 4072
rect 23155 3964 23520 3992
rect 23155 3961 23167 3964
rect 23109 3955 23167 3961
rect 19702 3924 19708 3936
rect 19536 3896 19708 3924
rect 18095 3893 18107 3896
rect 18049 3887 18107 3893
rect 19702 3884 19708 3896
rect 19760 3924 19766 3936
rect 20254 3924 20260 3936
rect 19760 3896 20260 3924
rect 19760 3884 19766 3896
rect 20254 3884 20260 3896
rect 20312 3884 20318 3936
rect 23382 3884 23388 3936
rect 23440 3884 23446 3936
rect 23658 3884 23664 3936
rect 23716 3884 23722 3936
rect 23750 3884 23756 3936
rect 23808 3884 23814 3936
rect 1104 3834 28888 3856
rect 1104 3782 4423 3834
rect 4475 3782 4487 3834
rect 4539 3782 4551 3834
rect 4603 3782 4615 3834
rect 4667 3782 4679 3834
rect 4731 3782 11369 3834
rect 11421 3782 11433 3834
rect 11485 3782 11497 3834
rect 11549 3782 11561 3834
rect 11613 3782 11625 3834
rect 11677 3782 18315 3834
rect 18367 3782 18379 3834
rect 18431 3782 18443 3834
rect 18495 3782 18507 3834
rect 18559 3782 18571 3834
rect 18623 3782 25261 3834
rect 25313 3782 25325 3834
rect 25377 3782 25389 3834
rect 25441 3782 25453 3834
rect 25505 3782 25517 3834
rect 25569 3782 28888 3834
rect 1104 3760 28888 3782
rect 18325 3723 18383 3729
rect 18325 3689 18337 3723
rect 18371 3720 18383 3723
rect 19426 3720 19432 3732
rect 18371 3692 19432 3720
rect 18371 3689 18383 3692
rect 18325 3683 18383 3689
rect 19426 3680 19432 3692
rect 19484 3680 19490 3732
rect 21450 3720 21456 3732
rect 20548 3692 21456 3720
rect 16574 3544 16580 3596
rect 16632 3584 16638 3596
rect 16632 3556 17908 3584
rect 16632 3544 16638 3556
rect 17880 3528 17908 3556
rect 19610 3544 19616 3596
rect 19668 3584 19674 3596
rect 19886 3584 19892 3596
rect 19668 3556 19892 3584
rect 19668 3544 19674 3556
rect 19886 3544 19892 3556
rect 19944 3544 19950 3596
rect 20165 3587 20223 3593
rect 20165 3553 20177 3587
rect 20211 3584 20223 3587
rect 20548 3584 20576 3692
rect 21450 3680 21456 3692
rect 21508 3680 21514 3732
rect 22186 3720 22192 3732
rect 22066 3692 22192 3720
rect 22066 3652 22094 3692
rect 22186 3680 22192 3692
rect 22244 3680 22250 3732
rect 22738 3680 22744 3732
rect 22796 3720 22802 3732
rect 23014 3720 23020 3732
rect 22796 3692 23020 3720
rect 22796 3680 22802 3692
rect 23014 3680 23020 3692
rect 23072 3720 23078 3732
rect 23109 3723 23167 3729
rect 23109 3720 23121 3723
rect 23072 3692 23121 3720
rect 23072 3680 23078 3692
rect 23109 3689 23121 3692
rect 23155 3720 23167 3723
rect 23382 3720 23388 3732
rect 23155 3692 23388 3720
rect 23155 3689 23167 3692
rect 23109 3683 23167 3689
rect 23382 3680 23388 3692
rect 23440 3680 23446 3732
rect 26142 3680 26148 3732
rect 26200 3680 26206 3732
rect 20211 3556 20576 3584
rect 20640 3624 22094 3652
rect 23569 3655 23627 3661
rect 20211 3553 20223 3556
rect 20165 3547 20223 3553
rect 17862 3476 17868 3528
rect 17920 3476 17926 3528
rect 17954 3476 17960 3528
rect 18012 3516 18018 3528
rect 18598 3516 18604 3528
rect 18012 3488 18604 3516
rect 18012 3476 18018 3488
rect 18598 3476 18604 3488
rect 18656 3516 18662 3528
rect 18877 3519 18935 3525
rect 18877 3516 18889 3519
rect 18656 3488 18889 3516
rect 18656 3476 18662 3488
rect 18877 3485 18889 3488
rect 18923 3485 18935 3519
rect 18877 3479 18935 3485
rect 20254 3476 20260 3528
rect 20312 3476 20318 3528
rect 20349 3519 20407 3525
rect 20349 3485 20361 3519
rect 20395 3516 20407 3519
rect 20640 3516 20668 3624
rect 23569 3621 23581 3655
rect 23615 3652 23627 3655
rect 23615 3624 24532 3652
rect 23615 3621 23627 3624
rect 23569 3615 23627 3621
rect 22557 3587 22615 3593
rect 22557 3584 22569 3587
rect 22066 3556 22569 3584
rect 20395 3488 20668 3516
rect 20395 3485 20407 3488
rect 20349 3479 20407 3485
rect 20806 3476 20812 3528
rect 20864 3476 20870 3528
rect 16850 3408 16856 3460
rect 16908 3408 16914 3460
rect 18509 3451 18567 3457
rect 18509 3417 18521 3451
rect 18555 3417 18567 3451
rect 20898 3448 20904 3460
rect 18509 3411 18567 3417
rect 18892 3420 20904 3448
rect 18524 3380 18552 3411
rect 18892 3392 18920 3420
rect 20898 3408 20904 3420
rect 20956 3408 20962 3460
rect 18874 3380 18880 3392
rect 18524 3352 18880 3380
rect 18874 3340 18880 3352
rect 18932 3340 18938 3392
rect 19245 3383 19303 3389
rect 19245 3349 19257 3383
rect 19291 3380 19303 3383
rect 19334 3380 19340 3392
rect 19291 3352 19340 3380
rect 19291 3349 19303 3352
rect 19245 3343 19303 3349
rect 19334 3340 19340 3352
rect 19392 3340 19398 3392
rect 20714 3340 20720 3392
rect 20772 3340 20778 3392
rect 21818 3340 21824 3392
rect 21876 3380 21882 3392
rect 22066 3380 22094 3556
rect 22557 3553 22569 3556
rect 22603 3584 22615 3587
rect 24210 3584 24216 3596
rect 22603 3556 24216 3584
rect 22603 3553 22615 3556
rect 22557 3547 22615 3553
rect 24210 3544 24216 3556
rect 24268 3584 24274 3596
rect 24397 3587 24455 3593
rect 24397 3584 24409 3587
rect 24268 3556 24409 3584
rect 24268 3544 24274 3556
rect 24397 3553 24409 3556
rect 24443 3553 24455 3587
rect 24504 3584 24532 3624
rect 24673 3587 24731 3593
rect 24673 3584 24685 3587
rect 24504 3556 24685 3584
rect 24397 3547 24455 3553
rect 24673 3553 24685 3556
rect 24719 3553 24731 3587
rect 24673 3547 24731 3553
rect 22833 3519 22891 3525
rect 22833 3516 22845 3519
rect 22572 3488 22845 3516
rect 22572 3460 22600 3488
rect 22833 3485 22845 3488
rect 22879 3485 22891 3519
rect 22833 3479 22891 3485
rect 23201 3519 23259 3525
rect 23201 3485 23213 3519
rect 23247 3485 23259 3519
rect 23201 3479 23259 3485
rect 22554 3408 22560 3460
rect 22612 3408 22618 3460
rect 21876 3352 22094 3380
rect 21876 3340 21882 3352
rect 22646 3340 22652 3392
rect 22704 3340 22710 3392
rect 22848 3380 22876 3479
rect 23106 3408 23112 3460
rect 23164 3448 23170 3460
rect 23216 3448 23244 3479
rect 23290 3476 23296 3528
rect 23348 3476 23354 3528
rect 23385 3519 23443 3525
rect 23385 3485 23397 3519
rect 23431 3516 23443 3519
rect 23474 3516 23480 3528
rect 23431 3488 23480 3516
rect 23431 3485 23443 3488
rect 23385 3479 23443 3485
rect 23474 3476 23480 3488
rect 23532 3476 23538 3528
rect 23569 3519 23627 3525
rect 23569 3485 23581 3519
rect 23615 3516 23627 3519
rect 23750 3516 23756 3528
rect 23615 3488 23756 3516
rect 23615 3485 23627 3488
rect 23569 3479 23627 3485
rect 23750 3476 23756 3488
rect 23808 3476 23814 3528
rect 23164 3420 23244 3448
rect 23164 3408 23170 3420
rect 25130 3408 25136 3460
rect 25188 3408 25194 3460
rect 23290 3380 23296 3392
rect 22848 3352 23296 3380
rect 23290 3340 23296 3352
rect 23348 3340 23354 3392
rect 1104 3290 28888 3312
rect 1104 3238 5083 3290
rect 5135 3238 5147 3290
rect 5199 3238 5211 3290
rect 5263 3238 5275 3290
rect 5327 3238 5339 3290
rect 5391 3238 12029 3290
rect 12081 3238 12093 3290
rect 12145 3238 12157 3290
rect 12209 3238 12221 3290
rect 12273 3238 12285 3290
rect 12337 3238 18975 3290
rect 19027 3238 19039 3290
rect 19091 3238 19103 3290
rect 19155 3238 19167 3290
rect 19219 3238 19231 3290
rect 19283 3238 25921 3290
rect 25973 3238 25985 3290
rect 26037 3238 26049 3290
rect 26101 3238 26113 3290
rect 26165 3238 26177 3290
rect 26229 3238 28888 3290
rect 1104 3216 28888 3238
rect 16850 3136 16856 3188
rect 16908 3176 16914 3188
rect 17221 3179 17279 3185
rect 17221 3176 17233 3179
rect 16908 3148 17233 3176
rect 16908 3136 16914 3148
rect 17221 3145 17233 3148
rect 17267 3145 17279 3179
rect 17221 3139 17279 3145
rect 17402 3136 17408 3188
rect 17460 3136 17466 3188
rect 19518 3176 19524 3188
rect 18156 3148 19524 3176
rect 17420 3049 17448 3136
rect 18156 3117 18184 3148
rect 19518 3136 19524 3148
rect 19576 3136 19582 3188
rect 19610 3136 19616 3188
rect 19668 3136 19674 3188
rect 19794 3176 19800 3188
rect 19720 3148 19800 3176
rect 18141 3111 18199 3117
rect 18141 3077 18153 3111
rect 18187 3077 18199 3111
rect 18141 3071 18199 3077
rect 18598 3068 18604 3120
rect 18656 3068 18662 3120
rect 17405 3043 17463 3049
rect 17405 3009 17417 3043
rect 17451 3009 17463 3043
rect 17405 3003 17463 3009
rect 17862 3000 17868 3052
rect 17920 3000 17926 3052
rect 19720 3049 19748 3148
rect 19794 3136 19800 3148
rect 19852 3176 19858 3188
rect 19852 3148 21864 3176
rect 19852 3136 19858 3148
rect 21726 3108 21732 3120
rect 21206 3094 21732 3108
rect 21192 3080 21732 3094
rect 19705 3043 19763 3049
rect 19705 3009 19717 3043
rect 19751 3009 19763 3043
rect 19705 3003 19763 3009
rect 21192 2984 21220 3080
rect 21726 3068 21732 3080
rect 21784 3068 21790 3120
rect 19978 2932 19984 2984
rect 20036 2932 20042 2984
rect 21174 2932 21180 2984
rect 21232 2932 21238 2984
rect 21450 2864 21456 2916
rect 21508 2864 21514 2916
rect 21744 2836 21772 3068
rect 21836 3052 21864 3148
rect 21818 3000 21824 3052
rect 21876 3000 21882 3052
rect 25130 3040 25136 3052
rect 23230 3026 25136 3040
rect 23216 3012 25136 3026
rect 22094 2932 22100 2984
rect 22152 2932 22158 2984
rect 23216 2836 23244 3012
rect 25130 3000 25136 3012
rect 25188 3000 25194 3052
rect 23474 2932 23480 2984
rect 23532 2972 23538 2984
rect 23569 2975 23627 2981
rect 23569 2972 23581 2975
rect 23532 2944 23581 2972
rect 23532 2932 23538 2944
rect 23569 2941 23581 2944
rect 23615 2972 23627 2975
rect 24213 2975 24271 2981
rect 24213 2972 24225 2975
rect 23615 2944 24225 2972
rect 23615 2941 23627 2944
rect 23569 2935 23627 2941
rect 24213 2941 24225 2944
rect 24259 2941 24271 2975
rect 24213 2935 24271 2941
rect 21744 2808 23244 2836
rect 23658 2796 23664 2848
rect 23716 2796 23722 2848
rect 1104 2746 28888 2768
rect 1104 2694 4423 2746
rect 4475 2694 4487 2746
rect 4539 2694 4551 2746
rect 4603 2694 4615 2746
rect 4667 2694 4679 2746
rect 4731 2694 11369 2746
rect 11421 2694 11433 2746
rect 11485 2694 11497 2746
rect 11549 2694 11561 2746
rect 11613 2694 11625 2746
rect 11677 2694 18315 2746
rect 18367 2694 18379 2746
rect 18431 2694 18443 2746
rect 18495 2694 18507 2746
rect 18559 2694 18571 2746
rect 18623 2694 25261 2746
rect 25313 2694 25325 2746
rect 25377 2694 25389 2746
rect 25441 2694 25453 2746
rect 25505 2694 25517 2746
rect 25569 2694 28888 2746
rect 1104 2672 28888 2694
rect 18138 2592 18144 2644
rect 18196 2592 18202 2644
rect 19978 2592 19984 2644
rect 20036 2632 20042 2644
rect 20257 2635 20315 2641
rect 20257 2632 20269 2635
rect 20036 2604 20269 2632
rect 20036 2592 20042 2604
rect 20257 2601 20269 2604
rect 20303 2601 20315 2635
rect 20257 2595 20315 2601
rect 21174 2592 21180 2644
rect 21232 2592 21238 2644
rect 21266 2592 21272 2644
rect 21324 2592 21330 2644
rect 22005 2635 22063 2641
rect 22005 2601 22017 2635
rect 22051 2632 22063 2635
rect 22094 2632 22100 2644
rect 22051 2604 22100 2632
rect 22051 2601 22063 2604
rect 22005 2595 22063 2601
rect 22094 2592 22100 2604
rect 22152 2592 22158 2644
rect 22741 2635 22799 2641
rect 22741 2601 22753 2635
rect 22787 2632 22799 2635
rect 23290 2632 23296 2644
rect 22787 2604 23296 2632
rect 22787 2601 22799 2604
rect 22741 2595 22799 2601
rect 23290 2592 23296 2604
rect 23348 2592 23354 2644
rect 19705 2567 19763 2573
rect 19705 2533 19717 2567
rect 19751 2564 19763 2567
rect 21284 2564 21312 2592
rect 23017 2567 23075 2573
rect 23017 2564 23029 2567
rect 19751 2536 21312 2564
rect 22204 2536 23029 2564
rect 19751 2533 19763 2536
rect 19705 2527 19763 2533
rect 1673 2499 1731 2505
rect 1673 2465 1685 2499
rect 1719 2496 1731 2499
rect 13538 2496 13544 2508
rect 1719 2468 13544 2496
rect 1719 2465 1731 2468
rect 1673 2459 1731 2465
rect 13538 2456 13544 2468
rect 13596 2456 13602 2508
rect 19334 2456 19340 2508
rect 19392 2456 19398 2508
rect 22204 2505 22232 2536
rect 23017 2533 23029 2536
rect 23063 2533 23075 2567
rect 23017 2527 23075 2533
rect 22189 2499 22247 2505
rect 22189 2465 22201 2499
rect 22235 2465 22247 2499
rect 22189 2459 22247 2465
rect 22646 2456 22652 2508
rect 22704 2456 22710 2508
rect 23032 2468 23428 2496
rect 14 2388 20 2440
rect 72 2428 78 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 72 2400 1409 2428
rect 72 2388 78 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 9122 2388 9128 2440
rect 9180 2388 9186 2440
rect 18046 2388 18052 2440
rect 18104 2428 18110 2440
rect 18325 2431 18383 2437
rect 18325 2428 18337 2431
rect 18104 2400 18337 2428
rect 18104 2388 18110 2400
rect 18325 2397 18337 2400
rect 18371 2397 18383 2431
rect 18325 2391 18383 2397
rect 19521 2431 19579 2437
rect 19521 2397 19533 2431
rect 19567 2428 19579 2431
rect 19610 2428 19616 2440
rect 19567 2400 19616 2428
rect 19567 2397 19579 2400
rect 19521 2391 19579 2397
rect 19610 2388 19616 2400
rect 19668 2388 19674 2440
rect 20441 2431 20499 2437
rect 20441 2397 20453 2431
rect 20487 2428 20499 2431
rect 20714 2428 20720 2440
rect 20487 2400 20720 2428
rect 20487 2397 20499 2400
rect 20441 2391 20499 2397
rect 20714 2388 20720 2400
rect 20772 2388 20778 2440
rect 20898 2388 20904 2440
rect 20956 2428 20962 2440
rect 23032 2437 23060 2468
rect 23400 2440 23428 2468
rect 23658 2456 23664 2508
rect 23716 2456 23722 2508
rect 21269 2431 21327 2437
rect 21269 2428 21281 2431
rect 20956 2400 21281 2428
rect 20956 2388 20962 2400
rect 21269 2397 21281 2400
rect 21315 2397 21327 2431
rect 21269 2391 21327 2397
rect 22281 2431 22339 2437
rect 22281 2397 22293 2431
rect 22327 2397 22339 2431
rect 22281 2391 22339 2397
rect 23017 2431 23075 2437
rect 23017 2397 23029 2431
rect 23063 2397 23075 2431
rect 23017 2391 23075 2397
rect 17126 2320 17132 2372
rect 17184 2360 17190 2372
rect 22296 2360 22324 2391
rect 23106 2388 23112 2440
rect 23164 2428 23170 2440
rect 23201 2431 23259 2437
rect 23201 2428 23213 2431
rect 23164 2400 23213 2428
rect 23164 2388 23170 2400
rect 23201 2397 23213 2400
rect 23247 2397 23259 2431
rect 23201 2391 23259 2397
rect 23382 2388 23388 2440
rect 23440 2388 23446 2440
rect 23676 2360 23704 2456
rect 27062 2388 27068 2440
rect 27120 2428 27126 2440
rect 27341 2431 27399 2437
rect 27341 2428 27353 2431
rect 27120 2400 27353 2428
rect 27120 2388 27126 2400
rect 27341 2397 27353 2400
rect 27387 2397 27399 2431
rect 27341 2391 27399 2397
rect 17184 2332 18920 2360
rect 22296 2332 23704 2360
rect 17184 2320 17190 2332
rect 9309 2295 9367 2301
rect 9309 2261 9321 2295
rect 9355 2292 9367 2295
rect 18782 2292 18788 2304
rect 9355 2264 18788 2292
rect 9355 2261 9367 2264
rect 9309 2255 9367 2261
rect 18782 2252 18788 2264
rect 18840 2252 18846 2304
rect 18892 2292 18920 2332
rect 27157 2295 27215 2301
rect 27157 2292 27169 2295
rect 18892 2264 27169 2292
rect 27157 2261 27169 2264
rect 27203 2261 27215 2295
rect 27157 2255 27215 2261
rect 1104 2202 28888 2224
rect 1104 2150 5083 2202
rect 5135 2150 5147 2202
rect 5199 2150 5211 2202
rect 5263 2150 5275 2202
rect 5327 2150 5339 2202
rect 5391 2150 12029 2202
rect 12081 2150 12093 2202
rect 12145 2150 12157 2202
rect 12209 2150 12221 2202
rect 12273 2150 12285 2202
rect 12337 2150 18975 2202
rect 19027 2150 19039 2202
rect 19091 2150 19103 2202
rect 19155 2150 19167 2202
rect 19219 2150 19231 2202
rect 19283 2150 25921 2202
rect 25973 2150 25985 2202
rect 26037 2150 26049 2202
rect 26101 2150 26113 2202
rect 26165 2150 26177 2202
rect 26229 2150 28888 2202
rect 1104 2128 28888 2150
<< via1 >>
rect 4423 27718 4475 27770
rect 4487 27718 4539 27770
rect 4551 27718 4603 27770
rect 4615 27718 4667 27770
rect 4679 27718 4731 27770
rect 11369 27718 11421 27770
rect 11433 27718 11485 27770
rect 11497 27718 11549 27770
rect 11561 27718 11613 27770
rect 11625 27718 11677 27770
rect 18315 27718 18367 27770
rect 18379 27718 18431 27770
rect 18443 27718 18495 27770
rect 18507 27718 18559 27770
rect 18571 27718 18623 27770
rect 25261 27718 25313 27770
rect 25325 27718 25377 27770
rect 25389 27718 25441 27770
rect 25453 27718 25505 27770
rect 25517 27718 25569 27770
rect 1492 27591 1544 27600
rect 1492 27557 1501 27591
rect 1501 27557 1535 27591
rect 1535 27557 1544 27591
rect 1492 27548 1544 27557
rect 7196 27548 7248 27600
rect 16120 27548 16172 27600
rect 21640 27548 21692 27600
rect 25136 27480 25188 27532
rect 17592 27412 17644 27464
rect 20996 27344 21048 27396
rect 15844 27276 15896 27328
rect 5083 27174 5135 27226
rect 5147 27174 5199 27226
rect 5211 27174 5263 27226
rect 5275 27174 5327 27226
rect 5339 27174 5391 27226
rect 12029 27174 12081 27226
rect 12093 27174 12145 27226
rect 12157 27174 12209 27226
rect 12221 27174 12273 27226
rect 12285 27174 12337 27226
rect 18975 27174 19027 27226
rect 19039 27174 19091 27226
rect 19103 27174 19155 27226
rect 19167 27174 19219 27226
rect 19231 27174 19283 27226
rect 25921 27174 25973 27226
rect 25985 27174 26037 27226
rect 26049 27174 26101 27226
rect 26113 27174 26165 27226
rect 26177 27174 26229 27226
rect 4423 26630 4475 26682
rect 4487 26630 4539 26682
rect 4551 26630 4603 26682
rect 4615 26630 4667 26682
rect 4679 26630 4731 26682
rect 11369 26630 11421 26682
rect 11433 26630 11485 26682
rect 11497 26630 11549 26682
rect 11561 26630 11613 26682
rect 11625 26630 11677 26682
rect 18315 26630 18367 26682
rect 18379 26630 18431 26682
rect 18443 26630 18495 26682
rect 18507 26630 18559 26682
rect 18571 26630 18623 26682
rect 25261 26630 25313 26682
rect 25325 26630 25377 26682
rect 25389 26630 25441 26682
rect 25453 26630 25505 26682
rect 25517 26630 25569 26682
rect 5083 26086 5135 26138
rect 5147 26086 5199 26138
rect 5211 26086 5263 26138
rect 5275 26086 5327 26138
rect 5339 26086 5391 26138
rect 12029 26086 12081 26138
rect 12093 26086 12145 26138
rect 12157 26086 12209 26138
rect 12221 26086 12273 26138
rect 12285 26086 12337 26138
rect 18975 26086 19027 26138
rect 19039 26086 19091 26138
rect 19103 26086 19155 26138
rect 19167 26086 19219 26138
rect 19231 26086 19283 26138
rect 25921 26086 25973 26138
rect 25985 26086 26037 26138
rect 26049 26086 26101 26138
rect 26113 26086 26165 26138
rect 26177 26086 26229 26138
rect 4423 25542 4475 25594
rect 4487 25542 4539 25594
rect 4551 25542 4603 25594
rect 4615 25542 4667 25594
rect 4679 25542 4731 25594
rect 11369 25542 11421 25594
rect 11433 25542 11485 25594
rect 11497 25542 11549 25594
rect 11561 25542 11613 25594
rect 11625 25542 11677 25594
rect 18315 25542 18367 25594
rect 18379 25542 18431 25594
rect 18443 25542 18495 25594
rect 18507 25542 18559 25594
rect 18571 25542 18623 25594
rect 25261 25542 25313 25594
rect 25325 25542 25377 25594
rect 25389 25542 25441 25594
rect 25453 25542 25505 25594
rect 25517 25542 25569 25594
rect 28264 25279 28316 25288
rect 28264 25245 28273 25279
rect 28273 25245 28307 25279
rect 28307 25245 28316 25279
rect 28264 25236 28316 25245
rect 28540 25279 28592 25288
rect 28540 25245 28549 25279
rect 28549 25245 28583 25279
rect 28583 25245 28592 25279
rect 28540 25236 28592 25245
rect 5083 24998 5135 25050
rect 5147 24998 5199 25050
rect 5211 24998 5263 25050
rect 5275 24998 5327 25050
rect 5339 24998 5391 25050
rect 12029 24998 12081 25050
rect 12093 24998 12145 25050
rect 12157 24998 12209 25050
rect 12221 24998 12273 25050
rect 12285 24998 12337 25050
rect 18975 24998 19027 25050
rect 19039 24998 19091 25050
rect 19103 24998 19155 25050
rect 19167 24998 19219 25050
rect 19231 24998 19283 25050
rect 25921 24998 25973 25050
rect 25985 24998 26037 25050
rect 26049 24998 26101 25050
rect 26113 24998 26165 25050
rect 26177 24998 26229 25050
rect 4423 24454 4475 24506
rect 4487 24454 4539 24506
rect 4551 24454 4603 24506
rect 4615 24454 4667 24506
rect 4679 24454 4731 24506
rect 11369 24454 11421 24506
rect 11433 24454 11485 24506
rect 11497 24454 11549 24506
rect 11561 24454 11613 24506
rect 11625 24454 11677 24506
rect 18315 24454 18367 24506
rect 18379 24454 18431 24506
rect 18443 24454 18495 24506
rect 18507 24454 18559 24506
rect 18571 24454 18623 24506
rect 25261 24454 25313 24506
rect 25325 24454 25377 24506
rect 25389 24454 25441 24506
rect 25453 24454 25505 24506
rect 25517 24454 25569 24506
rect 5083 23910 5135 23962
rect 5147 23910 5199 23962
rect 5211 23910 5263 23962
rect 5275 23910 5327 23962
rect 5339 23910 5391 23962
rect 12029 23910 12081 23962
rect 12093 23910 12145 23962
rect 12157 23910 12209 23962
rect 12221 23910 12273 23962
rect 12285 23910 12337 23962
rect 18975 23910 19027 23962
rect 19039 23910 19091 23962
rect 19103 23910 19155 23962
rect 19167 23910 19219 23962
rect 19231 23910 19283 23962
rect 25921 23910 25973 23962
rect 25985 23910 26037 23962
rect 26049 23910 26101 23962
rect 26113 23910 26165 23962
rect 26177 23910 26229 23962
rect 4423 23366 4475 23418
rect 4487 23366 4539 23418
rect 4551 23366 4603 23418
rect 4615 23366 4667 23418
rect 4679 23366 4731 23418
rect 11369 23366 11421 23418
rect 11433 23366 11485 23418
rect 11497 23366 11549 23418
rect 11561 23366 11613 23418
rect 11625 23366 11677 23418
rect 18315 23366 18367 23418
rect 18379 23366 18431 23418
rect 18443 23366 18495 23418
rect 18507 23366 18559 23418
rect 18571 23366 18623 23418
rect 25261 23366 25313 23418
rect 25325 23366 25377 23418
rect 25389 23366 25441 23418
rect 25453 23366 25505 23418
rect 25517 23366 25569 23418
rect 5083 22822 5135 22874
rect 5147 22822 5199 22874
rect 5211 22822 5263 22874
rect 5275 22822 5327 22874
rect 5339 22822 5391 22874
rect 12029 22822 12081 22874
rect 12093 22822 12145 22874
rect 12157 22822 12209 22874
rect 12221 22822 12273 22874
rect 12285 22822 12337 22874
rect 18975 22822 19027 22874
rect 19039 22822 19091 22874
rect 19103 22822 19155 22874
rect 19167 22822 19219 22874
rect 19231 22822 19283 22874
rect 25921 22822 25973 22874
rect 25985 22822 26037 22874
rect 26049 22822 26101 22874
rect 26113 22822 26165 22874
rect 26177 22822 26229 22874
rect 4423 22278 4475 22330
rect 4487 22278 4539 22330
rect 4551 22278 4603 22330
rect 4615 22278 4667 22330
rect 4679 22278 4731 22330
rect 11369 22278 11421 22330
rect 11433 22278 11485 22330
rect 11497 22278 11549 22330
rect 11561 22278 11613 22330
rect 11625 22278 11677 22330
rect 18315 22278 18367 22330
rect 18379 22278 18431 22330
rect 18443 22278 18495 22330
rect 18507 22278 18559 22330
rect 18571 22278 18623 22330
rect 25261 22278 25313 22330
rect 25325 22278 25377 22330
rect 25389 22278 25441 22330
rect 25453 22278 25505 22330
rect 25517 22278 25569 22330
rect 5083 21734 5135 21786
rect 5147 21734 5199 21786
rect 5211 21734 5263 21786
rect 5275 21734 5327 21786
rect 5339 21734 5391 21786
rect 12029 21734 12081 21786
rect 12093 21734 12145 21786
rect 12157 21734 12209 21786
rect 12221 21734 12273 21786
rect 12285 21734 12337 21786
rect 18975 21734 19027 21786
rect 19039 21734 19091 21786
rect 19103 21734 19155 21786
rect 19167 21734 19219 21786
rect 19231 21734 19283 21786
rect 25921 21734 25973 21786
rect 25985 21734 26037 21786
rect 26049 21734 26101 21786
rect 26113 21734 26165 21786
rect 26177 21734 26229 21786
rect 4423 21190 4475 21242
rect 4487 21190 4539 21242
rect 4551 21190 4603 21242
rect 4615 21190 4667 21242
rect 4679 21190 4731 21242
rect 11369 21190 11421 21242
rect 11433 21190 11485 21242
rect 11497 21190 11549 21242
rect 11561 21190 11613 21242
rect 11625 21190 11677 21242
rect 18315 21190 18367 21242
rect 18379 21190 18431 21242
rect 18443 21190 18495 21242
rect 18507 21190 18559 21242
rect 18571 21190 18623 21242
rect 25261 21190 25313 21242
rect 25325 21190 25377 21242
rect 25389 21190 25441 21242
rect 25453 21190 25505 21242
rect 25517 21190 25569 21242
rect 5083 20646 5135 20698
rect 5147 20646 5199 20698
rect 5211 20646 5263 20698
rect 5275 20646 5327 20698
rect 5339 20646 5391 20698
rect 12029 20646 12081 20698
rect 12093 20646 12145 20698
rect 12157 20646 12209 20698
rect 12221 20646 12273 20698
rect 12285 20646 12337 20698
rect 18975 20646 19027 20698
rect 19039 20646 19091 20698
rect 19103 20646 19155 20698
rect 19167 20646 19219 20698
rect 19231 20646 19283 20698
rect 25921 20646 25973 20698
rect 25985 20646 26037 20698
rect 26049 20646 26101 20698
rect 26113 20646 26165 20698
rect 26177 20646 26229 20698
rect 4423 20102 4475 20154
rect 4487 20102 4539 20154
rect 4551 20102 4603 20154
rect 4615 20102 4667 20154
rect 4679 20102 4731 20154
rect 11369 20102 11421 20154
rect 11433 20102 11485 20154
rect 11497 20102 11549 20154
rect 11561 20102 11613 20154
rect 11625 20102 11677 20154
rect 18315 20102 18367 20154
rect 18379 20102 18431 20154
rect 18443 20102 18495 20154
rect 18507 20102 18559 20154
rect 18571 20102 18623 20154
rect 25261 20102 25313 20154
rect 25325 20102 25377 20154
rect 25389 20102 25441 20154
rect 25453 20102 25505 20154
rect 25517 20102 25569 20154
rect 5083 19558 5135 19610
rect 5147 19558 5199 19610
rect 5211 19558 5263 19610
rect 5275 19558 5327 19610
rect 5339 19558 5391 19610
rect 12029 19558 12081 19610
rect 12093 19558 12145 19610
rect 12157 19558 12209 19610
rect 12221 19558 12273 19610
rect 12285 19558 12337 19610
rect 18975 19558 19027 19610
rect 19039 19558 19091 19610
rect 19103 19558 19155 19610
rect 19167 19558 19219 19610
rect 19231 19558 19283 19610
rect 25921 19558 25973 19610
rect 25985 19558 26037 19610
rect 26049 19558 26101 19610
rect 26113 19558 26165 19610
rect 26177 19558 26229 19610
rect 4423 19014 4475 19066
rect 4487 19014 4539 19066
rect 4551 19014 4603 19066
rect 4615 19014 4667 19066
rect 4679 19014 4731 19066
rect 11369 19014 11421 19066
rect 11433 19014 11485 19066
rect 11497 19014 11549 19066
rect 11561 19014 11613 19066
rect 11625 19014 11677 19066
rect 18315 19014 18367 19066
rect 18379 19014 18431 19066
rect 18443 19014 18495 19066
rect 18507 19014 18559 19066
rect 18571 19014 18623 19066
rect 25261 19014 25313 19066
rect 25325 19014 25377 19066
rect 25389 19014 25441 19066
rect 25453 19014 25505 19066
rect 25517 19014 25569 19066
rect 940 18708 992 18760
rect 13452 18708 13504 18760
rect 5083 18470 5135 18522
rect 5147 18470 5199 18522
rect 5211 18470 5263 18522
rect 5275 18470 5327 18522
rect 5339 18470 5391 18522
rect 12029 18470 12081 18522
rect 12093 18470 12145 18522
rect 12157 18470 12209 18522
rect 12221 18470 12273 18522
rect 12285 18470 12337 18522
rect 18975 18470 19027 18522
rect 19039 18470 19091 18522
rect 19103 18470 19155 18522
rect 19167 18470 19219 18522
rect 19231 18470 19283 18522
rect 25921 18470 25973 18522
rect 25985 18470 26037 18522
rect 26049 18470 26101 18522
rect 26113 18470 26165 18522
rect 26177 18470 26229 18522
rect 4423 17926 4475 17978
rect 4487 17926 4539 17978
rect 4551 17926 4603 17978
rect 4615 17926 4667 17978
rect 4679 17926 4731 17978
rect 11369 17926 11421 17978
rect 11433 17926 11485 17978
rect 11497 17926 11549 17978
rect 11561 17926 11613 17978
rect 11625 17926 11677 17978
rect 18315 17926 18367 17978
rect 18379 17926 18431 17978
rect 18443 17926 18495 17978
rect 18507 17926 18559 17978
rect 18571 17926 18623 17978
rect 25261 17926 25313 17978
rect 25325 17926 25377 17978
rect 25389 17926 25441 17978
rect 25453 17926 25505 17978
rect 25517 17926 25569 17978
rect 5083 17382 5135 17434
rect 5147 17382 5199 17434
rect 5211 17382 5263 17434
rect 5275 17382 5327 17434
rect 5339 17382 5391 17434
rect 12029 17382 12081 17434
rect 12093 17382 12145 17434
rect 12157 17382 12209 17434
rect 12221 17382 12273 17434
rect 12285 17382 12337 17434
rect 18975 17382 19027 17434
rect 19039 17382 19091 17434
rect 19103 17382 19155 17434
rect 19167 17382 19219 17434
rect 19231 17382 19283 17434
rect 25921 17382 25973 17434
rect 25985 17382 26037 17434
rect 26049 17382 26101 17434
rect 26113 17382 26165 17434
rect 26177 17382 26229 17434
rect 4423 16838 4475 16890
rect 4487 16838 4539 16890
rect 4551 16838 4603 16890
rect 4615 16838 4667 16890
rect 4679 16838 4731 16890
rect 11369 16838 11421 16890
rect 11433 16838 11485 16890
rect 11497 16838 11549 16890
rect 11561 16838 11613 16890
rect 11625 16838 11677 16890
rect 18315 16838 18367 16890
rect 18379 16838 18431 16890
rect 18443 16838 18495 16890
rect 18507 16838 18559 16890
rect 18571 16838 18623 16890
rect 25261 16838 25313 16890
rect 25325 16838 25377 16890
rect 25389 16838 25441 16890
rect 25453 16838 25505 16890
rect 25517 16838 25569 16890
rect 5083 16294 5135 16346
rect 5147 16294 5199 16346
rect 5211 16294 5263 16346
rect 5275 16294 5327 16346
rect 5339 16294 5391 16346
rect 12029 16294 12081 16346
rect 12093 16294 12145 16346
rect 12157 16294 12209 16346
rect 12221 16294 12273 16346
rect 12285 16294 12337 16346
rect 18975 16294 19027 16346
rect 19039 16294 19091 16346
rect 19103 16294 19155 16346
rect 19167 16294 19219 16346
rect 19231 16294 19283 16346
rect 25921 16294 25973 16346
rect 25985 16294 26037 16346
rect 26049 16294 26101 16346
rect 26113 16294 26165 16346
rect 26177 16294 26229 16346
rect 4423 15750 4475 15802
rect 4487 15750 4539 15802
rect 4551 15750 4603 15802
rect 4615 15750 4667 15802
rect 4679 15750 4731 15802
rect 11369 15750 11421 15802
rect 11433 15750 11485 15802
rect 11497 15750 11549 15802
rect 11561 15750 11613 15802
rect 11625 15750 11677 15802
rect 18315 15750 18367 15802
rect 18379 15750 18431 15802
rect 18443 15750 18495 15802
rect 18507 15750 18559 15802
rect 18571 15750 18623 15802
rect 25261 15750 25313 15802
rect 25325 15750 25377 15802
rect 25389 15750 25441 15802
rect 25453 15750 25505 15802
rect 25517 15750 25569 15802
rect 5083 15206 5135 15258
rect 5147 15206 5199 15258
rect 5211 15206 5263 15258
rect 5275 15206 5327 15258
rect 5339 15206 5391 15258
rect 12029 15206 12081 15258
rect 12093 15206 12145 15258
rect 12157 15206 12209 15258
rect 12221 15206 12273 15258
rect 12285 15206 12337 15258
rect 18975 15206 19027 15258
rect 19039 15206 19091 15258
rect 19103 15206 19155 15258
rect 19167 15206 19219 15258
rect 19231 15206 19283 15258
rect 25921 15206 25973 15258
rect 25985 15206 26037 15258
rect 26049 15206 26101 15258
rect 26113 15206 26165 15258
rect 26177 15206 26229 15258
rect 4423 14662 4475 14714
rect 4487 14662 4539 14714
rect 4551 14662 4603 14714
rect 4615 14662 4667 14714
rect 4679 14662 4731 14714
rect 11369 14662 11421 14714
rect 11433 14662 11485 14714
rect 11497 14662 11549 14714
rect 11561 14662 11613 14714
rect 11625 14662 11677 14714
rect 18315 14662 18367 14714
rect 18379 14662 18431 14714
rect 18443 14662 18495 14714
rect 18507 14662 18559 14714
rect 18571 14662 18623 14714
rect 25261 14662 25313 14714
rect 25325 14662 25377 14714
rect 25389 14662 25441 14714
rect 25453 14662 25505 14714
rect 25517 14662 25569 14714
rect 5083 14118 5135 14170
rect 5147 14118 5199 14170
rect 5211 14118 5263 14170
rect 5275 14118 5327 14170
rect 5339 14118 5391 14170
rect 12029 14118 12081 14170
rect 12093 14118 12145 14170
rect 12157 14118 12209 14170
rect 12221 14118 12273 14170
rect 12285 14118 12337 14170
rect 18975 14118 19027 14170
rect 19039 14118 19091 14170
rect 19103 14118 19155 14170
rect 19167 14118 19219 14170
rect 19231 14118 19283 14170
rect 25921 14118 25973 14170
rect 25985 14118 26037 14170
rect 26049 14118 26101 14170
rect 26113 14118 26165 14170
rect 26177 14118 26229 14170
rect 4423 13574 4475 13626
rect 4487 13574 4539 13626
rect 4551 13574 4603 13626
rect 4615 13574 4667 13626
rect 4679 13574 4731 13626
rect 11369 13574 11421 13626
rect 11433 13574 11485 13626
rect 11497 13574 11549 13626
rect 11561 13574 11613 13626
rect 11625 13574 11677 13626
rect 18315 13574 18367 13626
rect 18379 13574 18431 13626
rect 18443 13574 18495 13626
rect 18507 13574 18559 13626
rect 18571 13574 18623 13626
rect 25261 13574 25313 13626
rect 25325 13574 25377 13626
rect 25389 13574 25441 13626
rect 25453 13574 25505 13626
rect 25517 13574 25569 13626
rect 16672 13311 16724 13320
rect 16672 13277 16681 13311
rect 16681 13277 16715 13311
rect 16715 13277 16724 13311
rect 16672 13268 16724 13277
rect 16028 13175 16080 13184
rect 16028 13141 16037 13175
rect 16037 13141 16071 13175
rect 16071 13141 16080 13175
rect 16028 13132 16080 13141
rect 5083 13030 5135 13082
rect 5147 13030 5199 13082
rect 5211 13030 5263 13082
rect 5275 13030 5327 13082
rect 5339 13030 5391 13082
rect 12029 13030 12081 13082
rect 12093 13030 12145 13082
rect 12157 13030 12209 13082
rect 12221 13030 12273 13082
rect 12285 13030 12337 13082
rect 18975 13030 19027 13082
rect 19039 13030 19091 13082
rect 19103 13030 19155 13082
rect 19167 13030 19219 13082
rect 19231 13030 19283 13082
rect 25921 13030 25973 13082
rect 25985 13030 26037 13082
rect 26049 13030 26101 13082
rect 26113 13030 26165 13082
rect 26177 13030 26229 13082
rect 15844 12971 15896 12980
rect 15844 12937 15853 12971
rect 15853 12937 15887 12971
rect 15887 12937 15896 12971
rect 15844 12928 15896 12937
rect 16028 12928 16080 12980
rect 15476 12631 15528 12640
rect 15476 12597 15485 12631
rect 15485 12597 15519 12631
rect 15519 12597 15528 12631
rect 15476 12588 15528 12597
rect 16304 12631 16356 12640
rect 16304 12597 16313 12631
rect 16313 12597 16347 12631
rect 16347 12597 16356 12631
rect 16304 12588 16356 12597
rect 28264 12860 28316 12912
rect 19248 12835 19300 12844
rect 19248 12801 19257 12835
rect 19257 12801 19291 12835
rect 19291 12801 19300 12835
rect 19248 12792 19300 12801
rect 17316 12767 17368 12776
rect 17316 12733 17325 12767
rect 17325 12733 17359 12767
rect 17359 12733 17368 12767
rect 17316 12724 17368 12733
rect 17408 12724 17460 12776
rect 18880 12699 18932 12708
rect 18880 12665 18889 12699
rect 18889 12665 18923 12699
rect 18923 12665 18932 12699
rect 18880 12656 18932 12665
rect 17316 12588 17368 12640
rect 4423 12486 4475 12538
rect 4487 12486 4539 12538
rect 4551 12486 4603 12538
rect 4615 12486 4667 12538
rect 4679 12486 4731 12538
rect 11369 12486 11421 12538
rect 11433 12486 11485 12538
rect 11497 12486 11549 12538
rect 11561 12486 11613 12538
rect 11625 12486 11677 12538
rect 18315 12486 18367 12538
rect 18379 12486 18431 12538
rect 18443 12486 18495 12538
rect 18507 12486 18559 12538
rect 18571 12486 18623 12538
rect 25261 12486 25313 12538
rect 25325 12486 25377 12538
rect 25389 12486 25441 12538
rect 25453 12486 25505 12538
rect 25517 12486 25569 12538
rect 19248 12316 19300 12368
rect 16304 12248 16356 12300
rect 17960 12248 18012 12300
rect 15476 12180 15528 12232
rect 17592 12180 17644 12232
rect 16488 12112 16540 12164
rect 14924 12087 14976 12096
rect 14924 12053 14933 12087
rect 14933 12053 14967 12087
rect 14967 12053 14976 12087
rect 14924 12044 14976 12053
rect 15108 12044 15160 12096
rect 17408 12087 17460 12096
rect 17408 12053 17417 12087
rect 17417 12053 17451 12087
rect 17451 12053 17460 12087
rect 17408 12044 17460 12053
rect 5083 11942 5135 11994
rect 5147 11942 5199 11994
rect 5211 11942 5263 11994
rect 5275 11942 5327 11994
rect 5339 11942 5391 11994
rect 12029 11942 12081 11994
rect 12093 11942 12145 11994
rect 12157 11942 12209 11994
rect 12221 11942 12273 11994
rect 12285 11942 12337 11994
rect 18975 11942 19027 11994
rect 19039 11942 19091 11994
rect 19103 11942 19155 11994
rect 19167 11942 19219 11994
rect 19231 11942 19283 11994
rect 25921 11942 25973 11994
rect 25985 11942 26037 11994
rect 26049 11942 26101 11994
rect 26113 11942 26165 11994
rect 26177 11942 26229 11994
rect 14924 11840 14976 11892
rect 17592 11883 17644 11892
rect 17592 11849 17601 11883
rect 17601 11849 17635 11883
rect 17635 11849 17644 11883
rect 17592 11840 17644 11849
rect 21732 11772 21784 11824
rect 16488 11704 16540 11756
rect 18972 11747 19024 11756
rect 18972 11713 18981 11747
rect 18981 11713 19015 11747
rect 19015 11713 19024 11747
rect 18972 11704 19024 11713
rect 19248 11704 19300 11756
rect 14188 11500 14240 11552
rect 17316 11636 17368 11688
rect 17776 11679 17828 11688
rect 17776 11645 17785 11679
rect 17785 11645 17819 11679
rect 17819 11645 17828 11679
rect 17776 11636 17828 11645
rect 16672 11568 16724 11620
rect 18236 11568 18288 11620
rect 19984 11636 20036 11688
rect 20168 11679 20220 11688
rect 20168 11645 20177 11679
rect 20177 11645 20211 11679
rect 20211 11645 20220 11679
rect 20168 11636 20220 11645
rect 19340 11611 19392 11620
rect 19340 11577 19349 11611
rect 19349 11577 19383 11611
rect 19383 11577 19392 11611
rect 19340 11568 19392 11577
rect 15108 11500 15160 11552
rect 17224 11543 17276 11552
rect 17224 11509 17233 11543
rect 17233 11509 17267 11543
rect 17267 11509 17276 11543
rect 17224 11500 17276 11509
rect 17500 11500 17552 11552
rect 18052 11500 18104 11552
rect 19432 11543 19484 11552
rect 19432 11509 19441 11543
rect 19441 11509 19475 11543
rect 19475 11509 19484 11543
rect 19432 11500 19484 11509
rect 21640 11500 21692 11552
rect 4423 11398 4475 11450
rect 4487 11398 4539 11450
rect 4551 11398 4603 11450
rect 4615 11398 4667 11450
rect 4679 11398 4731 11450
rect 11369 11398 11421 11450
rect 11433 11398 11485 11450
rect 11497 11398 11549 11450
rect 11561 11398 11613 11450
rect 11625 11398 11677 11450
rect 18315 11398 18367 11450
rect 18379 11398 18431 11450
rect 18443 11398 18495 11450
rect 18507 11398 18559 11450
rect 18571 11398 18623 11450
rect 25261 11398 25313 11450
rect 25325 11398 25377 11450
rect 25389 11398 25441 11450
rect 25453 11398 25505 11450
rect 25517 11398 25569 11450
rect 16580 11296 16632 11348
rect 19248 11339 19300 11348
rect 19248 11305 19257 11339
rect 19257 11305 19291 11339
rect 19291 11305 19300 11339
rect 19248 11296 19300 11305
rect 20996 11339 21048 11348
rect 20996 11305 21005 11339
rect 21005 11305 21039 11339
rect 21039 11305 21048 11339
rect 20996 11296 21048 11305
rect 21456 11296 21508 11348
rect 18052 11228 18104 11280
rect 13452 11203 13504 11212
rect 13452 11169 13461 11203
rect 13461 11169 13495 11203
rect 13495 11169 13504 11203
rect 13452 11160 13504 11169
rect 13820 11160 13872 11212
rect 15016 11160 15068 11212
rect 13544 11135 13596 11144
rect 13544 11101 13553 11135
rect 13553 11101 13587 11135
rect 13587 11101 13596 11135
rect 13544 11092 13596 11101
rect 14188 11135 14240 11144
rect 14188 11101 14197 11135
rect 14197 11101 14231 11135
rect 14231 11101 14240 11135
rect 14188 11092 14240 11101
rect 16488 11160 16540 11212
rect 15752 11024 15804 11076
rect 17776 11160 17828 11212
rect 18788 11092 18840 11144
rect 19340 11092 19392 11144
rect 20720 11135 20772 11144
rect 20720 11101 20729 11135
rect 20729 11101 20763 11135
rect 20763 11101 20772 11135
rect 20720 11092 20772 11101
rect 15936 10999 15988 11008
rect 15936 10965 15945 10999
rect 15945 10965 15979 10999
rect 15979 10965 15988 10999
rect 15936 10956 15988 10965
rect 16304 10956 16356 11008
rect 17316 10956 17368 11008
rect 18144 10956 18196 11008
rect 22008 11024 22060 11076
rect 22468 11067 22520 11076
rect 22468 11033 22477 11067
rect 22477 11033 22511 11067
rect 22511 11033 22520 11067
rect 22468 11024 22520 11033
rect 18880 10956 18932 11008
rect 22560 10956 22612 11008
rect 5083 10854 5135 10906
rect 5147 10854 5199 10906
rect 5211 10854 5263 10906
rect 5275 10854 5327 10906
rect 5339 10854 5391 10906
rect 12029 10854 12081 10906
rect 12093 10854 12145 10906
rect 12157 10854 12209 10906
rect 12221 10854 12273 10906
rect 12285 10854 12337 10906
rect 18975 10854 19027 10906
rect 19039 10854 19091 10906
rect 19103 10854 19155 10906
rect 19167 10854 19219 10906
rect 19231 10854 19283 10906
rect 25921 10854 25973 10906
rect 25985 10854 26037 10906
rect 26049 10854 26101 10906
rect 26113 10854 26165 10906
rect 26177 10854 26229 10906
rect 13820 10752 13872 10804
rect 15016 10795 15068 10804
rect 15016 10761 15025 10795
rect 15025 10761 15059 10795
rect 15059 10761 15068 10795
rect 15016 10752 15068 10761
rect 17224 10752 17276 10804
rect 17316 10795 17368 10804
rect 17316 10761 17325 10795
rect 17325 10761 17359 10795
rect 17359 10761 17368 10795
rect 17316 10752 17368 10761
rect 18144 10752 18196 10804
rect 16396 10616 16448 10668
rect 17960 10659 18012 10668
rect 17960 10625 17969 10659
rect 17969 10625 18003 10659
rect 18003 10625 18012 10659
rect 17960 10616 18012 10625
rect 20720 10752 20772 10804
rect 22468 10752 22520 10804
rect 19708 10684 19760 10736
rect 23940 10752 23992 10804
rect 21272 10659 21324 10668
rect 21272 10625 21281 10659
rect 21281 10625 21315 10659
rect 21315 10625 21324 10659
rect 21272 10616 21324 10625
rect 21824 10616 21876 10668
rect 15936 10591 15988 10600
rect 15936 10557 15945 10591
rect 15945 10557 15979 10591
rect 15979 10557 15988 10591
rect 15936 10548 15988 10557
rect 16488 10548 16540 10600
rect 16580 10548 16632 10600
rect 17776 10591 17828 10600
rect 17776 10557 17785 10591
rect 17785 10557 17819 10591
rect 17819 10557 17828 10591
rect 17776 10548 17828 10557
rect 18236 10548 18288 10600
rect 19432 10548 19484 10600
rect 21916 10523 21968 10532
rect 21916 10489 21925 10523
rect 21925 10489 21959 10523
rect 21959 10489 21968 10523
rect 21916 10480 21968 10489
rect 15016 10412 15068 10464
rect 18236 10412 18288 10464
rect 18696 10412 18748 10464
rect 19984 10412 20036 10464
rect 21548 10412 21600 10464
rect 22284 10659 22336 10668
rect 22284 10625 22293 10659
rect 22293 10625 22327 10659
rect 22327 10625 22336 10659
rect 22284 10616 22336 10625
rect 24032 10616 24084 10668
rect 22560 10548 22612 10600
rect 24308 10412 24360 10464
rect 4423 10310 4475 10362
rect 4487 10310 4539 10362
rect 4551 10310 4603 10362
rect 4615 10310 4667 10362
rect 4679 10310 4731 10362
rect 11369 10310 11421 10362
rect 11433 10310 11485 10362
rect 11497 10310 11549 10362
rect 11561 10310 11613 10362
rect 11625 10310 11677 10362
rect 18315 10310 18367 10362
rect 18379 10310 18431 10362
rect 18443 10310 18495 10362
rect 18507 10310 18559 10362
rect 18571 10310 18623 10362
rect 25261 10310 25313 10362
rect 25325 10310 25377 10362
rect 25389 10310 25441 10362
rect 25453 10310 25505 10362
rect 25517 10310 25569 10362
rect 15108 10208 15160 10260
rect 16304 10208 16356 10260
rect 18696 10208 18748 10260
rect 18788 10208 18840 10260
rect 20812 10208 20864 10260
rect 22008 10208 22060 10260
rect 18236 10140 18288 10192
rect 15752 10004 15804 10056
rect 21364 10140 21416 10192
rect 20720 10072 20772 10124
rect 14372 9979 14424 9988
rect 14372 9945 14381 9979
rect 14381 9945 14415 9979
rect 14415 9945 14424 9979
rect 14372 9936 14424 9945
rect 21088 10047 21140 10056
rect 21088 10013 21097 10047
rect 21097 10013 21131 10047
rect 21131 10013 21140 10047
rect 21088 10004 21140 10013
rect 21180 10047 21232 10056
rect 21180 10013 21189 10047
rect 21189 10013 21223 10047
rect 21223 10013 21232 10047
rect 21180 10004 21232 10013
rect 21640 10072 21692 10124
rect 22560 10072 22612 10124
rect 23204 10072 23256 10124
rect 21824 10047 21876 10056
rect 21824 10013 21833 10047
rect 21833 10013 21867 10047
rect 21867 10013 21876 10047
rect 21824 10004 21876 10013
rect 22008 10047 22060 10056
rect 22008 10013 22017 10047
rect 22017 10013 22051 10047
rect 22051 10013 22060 10047
rect 22008 10004 22060 10013
rect 18696 9936 18748 9988
rect 18880 9936 18932 9988
rect 19616 9936 19668 9988
rect 20260 9979 20312 9988
rect 20260 9945 20269 9979
rect 20269 9945 20303 9979
rect 20303 9945 20312 9979
rect 20260 9936 20312 9945
rect 15936 9911 15988 9920
rect 15936 9877 15945 9911
rect 15945 9877 15979 9911
rect 15979 9877 15988 9911
rect 15936 9868 15988 9877
rect 17592 9868 17644 9920
rect 20536 9868 20588 9920
rect 20904 9911 20956 9920
rect 20904 9877 20913 9911
rect 20913 9877 20947 9911
rect 20947 9877 20956 9911
rect 20904 9868 20956 9877
rect 21548 9936 21600 9988
rect 22468 9979 22520 9988
rect 22468 9945 22477 9979
rect 22477 9945 22511 9979
rect 22511 9945 22520 9979
rect 22468 9936 22520 9945
rect 24032 9936 24084 9988
rect 24308 9936 24360 9988
rect 22560 9868 22612 9920
rect 5083 9766 5135 9818
rect 5147 9766 5199 9818
rect 5211 9766 5263 9818
rect 5275 9766 5327 9818
rect 5339 9766 5391 9818
rect 12029 9766 12081 9818
rect 12093 9766 12145 9818
rect 12157 9766 12209 9818
rect 12221 9766 12273 9818
rect 12285 9766 12337 9818
rect 18975 9766 19027 9818
rect 19039 9766 19091 9818
rect 19103 9766 19155 9818
rect 19167 9766 19219 9818
rect 19231 9766 19283 9818
rect 25921 9766 25973 9818
rect 25985 9766 26037 9818
rect 26049 9766 26101 9818
rect 26113 9766 26165 9818
rect 26177 9766 26229 9818
rect 14372 9664 14424 9716
rect 15936 9664 15988 9716
rect 19616 9707 19668 9716
rect 19616 9673 19625 9707
rect 19625 9673 19659 9707
rect 19659 9673 19668 9707
rect 19616 9664 19668 9673
rect 20812 9664 20864 9716
rect 21916 9664 21968 9716
rect 22284 9664 22336 9716
rect 22468 9664 22520 9716
rect 13544 9528 13596 9580
rect 14740 9460 14792 9512
rect 14740 9324 14792 9376
rect 17408 9571 17460 9580
rect 17408 9537 17417 9571
rect 17417 9537 17451 9571
rect 17451 9537 17460 9571
rect 17408 9528 17460 9537
rect 18236 9528 18288 9580
rect 18788 9528 18840 9580
rect 16396 9460 16448 9512
rect 16488 9460 16540 9512
rect 17684 9503 17736 9512
rect 17684 9469 17693 9503
rect 17693 9469 17727 9503
rect 17727 9469 17736 9503
rect 17684 9460 17736 9469
rect 16764 9367 16816 9376
rect 16764 9333 16773 9367
rect 16773 9333 16807 9367
rect 16807 9333 16816 9367
rect 16764 9324 16816 9333
rect 17224 9324 17276 9376
rect 17316 9324 17368 9376
rect 17684 9324 17736 9376
rect 18144 9392 18196 9444
rect 18788 9392 18840 9444
rect 20904 9528 20956 9580
rect 20996 9571 21048 9580
rect 20996 9537 21005 9571
rect 21005 9537 21039 9571
rect 21039 9537 21048 9571
rect 20996 9528 21048 9537
rect 21364 9596 21416 9648
rect 22008 9596 22060 9648
rect 21640 9528 21692 9580
rect 19432 9392 19484 9444
rect 20076 9503 20128 9512
rect 20076 9469 20085 9503
rect 20085 9469 20119 9503
rect 20119 9469 20128 9503
rect 20076 9460 20128 9469
rect 20536 9503 20588 9512
rect 20536 9469 20545 9503
rect 20545 9469 20579 9503
rect 20579 9469 20588 9503
rect 20536 9460 20588 9469
rect 20168 9392 20220 9444
rect 21088 9392 21140 9444
rect 22652 9503 22704 9512
rect 22652 9469 22661 9503
rect 22661 9469 22695 9503
rect 22695 9469 22704 9503
rect 22652 9460 22704 9469
rect 18236 9324 18288 9376
rect 19248 9367 19300 9376
rect 19248 9333 19257 9367
rect 19257 9333 19291 9367
rect 19291 9333 19300 9367
rect 19248 9324 19300 9333
rect 19340 9324 19392 9376
rect 20812 9324 20864 9376
rect 20996 9324 21048 9376
rect 21180 9324 21232 9376
rect 22284 9324 22336 9376
rect 23388 9392 23440 9444
rect 24124 9460 24176 9512
rect 4423 9222 4475 9274
rect 4487 9222 4539 9274
rect 4551 9222 4603 9274
rect 4615 9222 4667 9274
rect 4679 9222 4731 9274
rect 11369 9222 11421 9274
rect 11433 9222 11485 9274
rect 11497 9222 11549 9274
rect 11561 9222 11613 9274
rect 11625 9222 11677 9274
rect 18315 9222 18367 9274
rect 18379 9222 18431 9274
rect 18443 9222 18495 9274
rect 18507 9222 18559 9274
rect 18571 9222 18623 9274
rect 25261 9222 25313 9274
rect 25325 9222 25377 9274
rect 25389 9222 25441 9274
rect 25453 9222 25505 9274
rect 25517 9222 25569 9274
rect 940 8916 992 8968
rect 15016 9027 15068 9036
rect 15016 8993 15025 9027
rect 15025 8993 15059 9027
rect 15059 8993 15068 9027
rect 17776 9120 17828 9172
rect 19248 9120 19300 9172
rect 20260 9120 20312 9172
rect 20720 9120 20772 9172
rect 21272 9120 21324 9172
rect 17040 9052 17092 9104
rect 15016 8984 15068 8993
rect 15936 9027 15988 9036
rect 15936 8993 15945 9027
rect 15945 8993 15979 9027
rect 15979 8993 15988 9027
rect 15936 8984 15988 8993
rect 17132 9027 17184 9036
rect 17132 8993 17141 9027
rect 17141 8993 17175 9027
rect 17175 8993 17184 9027
rect 17132 8984 17184 8993
rect 17500 9027 17552 9036
rect 17500 8993 17534 9027
rect 17534 8993 17552 9027
rect 17500 8984 17552 8993
rect 17684 9027 17736 9036
rect 17684 8993 17693 9027
rect 17693 8993 17727 9027
rect 17727 8993 17736 9027
rect 19432 9052 19484 9104
rect 20812 9052 20864 9104
rect 22008 9052 22060 9104
rect 22284 9163 22336 9172
rect 22284 9129 22293 9163
rect 22293 9129 22327 9163
rect 22327 9129 22336 9163
rect 22284 9120 22336 9129
rect 17684 8984 17736 8993
rect 16028 8959 16080 8968
rect 16028 8925 16037 8959
rect 16037 8925 16071 8959
rect 16071 8925 16080 8959
rect 16028 8916 16080 8925
rect 16396 8916 16448 8968
rect 18880 8984 18932 9036
rect 18604 8959 18656 8968
rect 18604 8925 18613 8959
rect 18613 8925 18647 8959
rect 18647 8925 18656 8959
rect 18604 8916 18656 8925
rect 20904 8984 20956 9036
rect 14740 8891 14792 8900
rect 14740 8857 14749 8891
rect 14749 8857 14783 8891
rect 14783 8857 14792 8891
rect 14740 8848 14792 8857
rect 20996 8959 21048 8968
rect 20996 8925 21005 8959
rect 21005 8925 21039 8959
rect 21039 8925 21048 8959
rect 20996 8916 21048 8925
rect 21364 8916 21416 8968
rect 21456 8959 21508 8968
rect 21456 8925 21465 8959
rect 21465 8925 21499 8959
rect 21499 8925 21508 8959
rect 21456 8916 21508 8925
rect 21824 8916 21876 8968
rect 22652 8916 22704 8968
rect 14096 8823 14148 8832
rect 14096 8789 14105 8823
rect 14105 8789 14139 8823
rect 14139 8789 14148 8823
rect 14096 8780 14148 8789
rect 16212 8823 16264 8832
rect 16212 8789 16221 8823
rect 16221 8789 16255 8823
rect 16255 8789 16264 8823
rect 16212 8780 16264 8789
rect 18236 8780 18288 8832
rect 19340 8780 19392 8832
rect 20352 8780 20404 8832
rect 20536 8780 20588 8832
rect 21456 8780 21508 8832
rect 21548 8823 21600 8832
rect 21548 8789 21557 8823
rect 21557 8789 21591 8823
rect 21591 8789 21600 8823
rect 21548 8780 21600 8789
rect 22468 8780 22520 8832
rect 22652 8823 22704 8832
rect 22652 8789 22661 8823
rect 22661 8789 22695 8823
rect 22695 8789 22704 8823
rect 22652 8780 22704 8789
rect 22836 8891 22888 8900
rect 22836 8857 22870 8891
rect 22870 8857 22888 8891
rect 23388 8916 23440 8968
rect 24768 8916 24820 8968
rect 22836 8848 22888 8857
rect 23480 8780 23532 8832
rect 23756 8823 23808 8832
rect 23756 8789 23765 8823
rect 23765 8789 23799 8823
rect 23799 8789 23808 8823
rect 23756 8780 23808 8789
rect 24124 8780 24176 8832
rect 5083 8678 5135 8730
rect 5147 8678 5199 8730
rect 5211 8678 5263 8730
rect 5275 8678 5327 8730
rect 5339 8678 5391 8730
rect 12029 8678 12081 8730
rect 12093 8678 12145 8730
rect 12157 8678 12209 8730
rect 12221 8678 12273 8730
rect 12285 8678 12337 8730
rect 18975 8678 19027 8730
rect 19039 8678 19091 8730
rect 19103 8678 19155 8730
rect 19167 8678 19219 8730
rect 19231 8678 19283 8730
rect 25921 8678 25973 8730
rect 25985 8678 26037 8730
rect 26049 8678 26101 8730
rect 26113 8678 26165 8730
rect 26177 8678 26229 8730
rect 15108 8576 15160 8628
rect 15936 8576 15988 8628
rect 16028 8576 16080 8628
rect 14096 8508 14148 8560
rect 15752 8508 15804 8560
rect 19340 8576 19392 8628
rect 20352 8576 20404 8628
rect 20812 8576 20864 8628
rect 17224 8508 17276 8560
rect 18144 8508 18196 8560
rect 18696 8508 18748 8560
rect 16396 8372 16448 8424
rect 17776 8440 17828 8492
rect 19984 8483 20036 8492
rect 19984 8449 19993 8483
rect 19993 8449 20027 8483
rect 20027 8449 20036 8483
rect 19984 8440 20036 8449
rect 20260 8483 20312 8492
rect 20260 8449 20269 8483
rect 20269 8449 20303 8483
rect 20303 8449 20312 8483
rect 20260 8440 20312 8449
rect 21548 8576 21600 8628
rect 22008 8576 22060 8628
rect 22652 8576 22704 8628
rect 23388 8576 23440 8628
rect 21088 8440 21140 8492
rect 21456 8440 21508 8492
rect 20168 8372 20220 8424
rect 20536 8415 20588 8424
rect 20536 8381 20545 8415
rect 20545 8381 20579 8415
rect 20579 8381 20588 8415
rect 20536 8372 20588 8381
rect 21180 8415 21232 8424
rect 21180 8381 21189 8415
rect 21189 8381 21223 8415
rect 21223 8381 21232 8415
rect 21180 8372 21232 8381
rect 21640 8483 21692 8492
rect 21640 8449 21649 8483
rect 21649 8449 21683 8483
rect 21683 8449 21692 8483
rect 21640 8440 21692 8449
rect 23480 8508 23532 8560
rect 23756 8576 23808 8628
rect 24032 8508 24084 8560
rect 22560 8440 22612 8492
rect 23204 8372 23256 8424
rect 24216 8236 24268 8288
rect 24768 8236 24820 8288
rect 4423 8134 4475 8186
rect 4487 8134 4539 8186
rect 4551 8134 4603 8186
rect 4615 8134 4667 8186
rect 4679 8134 4731 8186
rect 11369 8134 11421 8186
rect 11433 8134 11485 8186
rect 11497 8134 11549 8186
rect 11561 8134 11613 8186
rect 11625 8134 11677 8186
rect 18315 8134 18367 8186
rect 18379 8134 18431 8186
rect 18443 8134 18495 8186
rect 18507 8134 18559 8186
rect 18571 8134 18623 8186
rect 25261 8134 25313 8186
rect 25325 8134 25377 8186
rect 25389 8134 25441 8186
rect 25453 8134 25505 8186
rect 25517 8134 25569 8186
rect 15108 8032 15160 8084
rect 17132 8032 17184 8084
rect 17500 8032 17552 8084
rect 18696 8032 18748 8084
rect 17868 7964 17920 8016
rect 18328 7964 18380 8016
rect 20260 8032 20312 8084
rect 21180 8032 21232 8084
rect 22836 8032 22888 8084
rect 23480 8032 23532 8084
rect 23940 8075 23992 8084
rect 23940 8041 23949 8075
rect 23949 8041 23983 8075
rect 23983 8041 23992 8075
rect 23940 8032 23992 8041
rect 24768 8032 24820 8084
rect 20720 7964 20772 8016
rect 20812 7964 20864 8016
rect 17684 7871 17736 7880
rect 17684 7837 17693 7871
rect 17693 7837 17727 7871
rect 17727 7837 17736 7871
rect 17684 7828 17736 7837
rect 17776 7871 17828 7880
rect 17776 7837 17785 7871
rect 17785 7837 17819 7871
rect 17819 7837 17828 7871
rect 17776 7828 17828 7837
rect 18236 7828 18288 7880
rect 18696 7871 18748 7880
rect 18696 7837 18705 7871
rect 18705 7837 18739 7871
rect 18739 7837 18748 7871
rect 18696 7828 18748 7837
rect 19432 7828 19484 7880
rect 20996 7896 21048 7948
rect 20076 7828 20128 7880
rect 20168 7760 20220 7812
rect 20444 7760 20496 7812
rect 17040 7692 17092 7744
rect 18236 7692 18288 7744
rect 20904 7828 20956 7880
rect 21824 7871 21876 7880
rect 21824 7837 21833 7871
rect 21833 7837 21867 7871
rect 21867 7837 21876 7871
rect 21824 7828 21876 7837
rect 22468 7964 22520 8016
rect 24032 7896 24084 7948
rect 24124 7939 24176 7948
rect 24124 7905 24133 7939
rect 24133 7905 24167 7939
rect 24167 7905 24176 7939
rect 24124 7896 24176 7905
rect 20720 7692 20772 7744
rect 22560 7692 22612 7744
rect 23204 7735 23256 7744
rect 23204 7701 23213 7735
rect 23213 7701 23247 7735
rect 23247 7701 23256 7735
rect 23204 7692 23256 7701
rect 24216 7803 24268 7812
rect 24216 7769 24225 7803
rect 24225 7769 24259 7803
rect 24259 7769 24268 7803
rect 24216 7760 24268 7769
rect 24308 7692 24360 7744
rect 28264 7760 28316 7812
rect 24860 7735 24912 7744
rect 24860 7701 24869 7735
rect 24869 7701 24903 7735
rect 24903 7701 24912 7735
rect 24860 7692 24912 7701
rect 25044 7692 25096 7744
rect 5083 7590 5135 7642
rect 5147 7590 5199 7642
rect 5211 7590 5263 7642
rect 5275 7590 5327 7642
rect 5339 7590 5391 7642
rect 12029 7590 12081 7642
rect 12093 7590 12145 7642
rect 12157 7590 12209 7642
rect 12221 7590 12273 7642
rect 12285 7590 12337 7642
rect 18975 7590 19027 7642
rect 19039 7590 19091 7642
rect 19103 7590 19155 7642
rect 19167 7590 19219 7642
rect 19231 7590 19283 7642
rect 25921 7590 25973 7642
rect 25985 7590 26037 7642
rect 26049 7590 26101 7642
rect 26113 7590 26165 7642
rect 26177 7590 26229 7642
rect 16396 7488 16448 7540
rect 15752 7420 15804 7472
rect 16212 7463 16264 7472
rect 16212 7429 16221 7463
rect 16221 7429 16255 7463
rect 16255 7429 16264 7463
rect 16212 7420 16264 7429
rect 17500 7488 17552 7540
rect 17684 7488 17736 7540
rect 18328 7531 18380 7540
rect 18328 7497 18337 7531
rect 18337 7497 18371 7531
rect 18371 7497 18380 7531
rect 18328 7488 18380 7497
rect 18696 7488 18748 7540
rect 20720 7531 20772 7540
rect 20720 7497 20747 7531
rect 20747 7497 20772 7531
rect 20720 7488 20772 7497
rect 20996 7488 21048 7540
rect 22468 7531 22520 7540
rect 22468 7497 22477 7531
rect 22477 7497 22511 7531
rect 22511 7497 22520 7531
rect 22468 7488 22520 7497
rect 19708 7420 19760 7472
rect 20444 7463 20496 7472
rect 20444 7429 20453 7463
rect 20453 7429 20487 7463
rect 20487 7429 20496 7463
rect 20444 7420 20496 7429
rect 17592 7352 17644 7404
rect 21456 7463 21508 7472
rect 21456 7429 21465 7463
rect 21465 7429 21499 7463
rect 21499 7429 21508 7463
rect 21456 7420 21508 7429
rect 21180 7395 21232 7404
rect 21180 7361 21189 7395
rect 21189 7361 21223 7395
rect 21223 7361 21232 7395
rect 21180 7352 21232 7361
rect 21640 7395 21692 7404
rect 21640 7361 21649 7395
rect 21649 7361 21683 7395
rect 21683 7361 21692 7395
rect 21640 7352 21692 7361
rect 16580 7284 16632 7336
rect 18696 7327 18748 7336
rect 18696 7293 18705 7327
rect 18705 7293 18739 7327
rect 18739 7293 18748 7327
rect 18696 7284 18748 7293
rect 21916 7395 21968 7404
rect 21916 7361 21925 7395
rect 21925 7361 21959 7395
rect 21959 7361 21968 7395
rect 21916 7352 21968 7361
rect 22192 7395 22244 7404
rect 22192 7361 22201 7395
rect 22201 7361 22235 7395
rect 22235 7361 22244 7395
rect 22192 7352 22244 7361
rect 20904 7216 20956 7268
rect 21180 7148 21232 7200
rect 22376 7284 22428 7336
rect 22560 7327 22612 7336
rect 22560 7293 22569 7327
rect 22569 7293 22603 7327
rect 22603 7293 22612 7327
rect 22560 7284 22612 7293
rect 22744 7327 22796 7336
rect 22744 7293 22753 7327
rect 22753 7293 22787 7327
rect 22787 7293 22796 7327
rect 22744 7284 22796 7293
rect 22836 7327 22888 7336
rect 22836 7293 22845 7327
rect 22845 7293 22879 7327
rect 22879 7293 22888 7327
rect 22836 7284 22888 7293
rect 23020 7327 23072 7336
rect 23020 7293 23029 7327
rect 23029 7293 23063 7327
rect 23063 7293 23072 7327
rect 23020 7284 23072 7293
rect 23204 7284 23256 7336
rect 23664 7327 23716 7336
rect 23664 7293 23673 7327
rect 23673 7293 23707 7327
rect 23707 7293 23716 7327
rect 23664 7284 23716 7293
rect 22560 7148 22612 7200
rect 24860 7216 24912 7268
rect 24952 7148 25004 7200
rect 4423 7046 4475 7098
rect 4487 7046 4539 7098
rect 4551 7046 4603 7098
rect 4615 7046 4667 7098
rect 4679 7046 4731 7098
rect 11369 7046 11421 7098
rect 11433 7046 11485 7098
rect 11497 7046 11549 7098
rect 11561 7046 11613 7098
rect 11625 7046 11677 7098
rect 18315 7046 18367 7098
rect 18379 7046 18431 7098
rect 18443 7046 18495 7098
rect 18507 7046 18559 7098
rect 18571 7046 18623 7098
rect 25261 7046 25313 7098
rect 25325 7046 25377 7098
rect 25389 7046 25441 7098
rect 25453 7046 25505 7098
rect 25517 7046 25569 7098
rect 17040 6944 17092 6996
rect 17684 6944 17736 6996
rect 18696 6987 18748 6996
rect 18696 6953 18705 6987
rect 18705 6953 18739 6987
rect 18739 6953 18748 6987
rect 18696 6944 18748 6953
rect 23664 6944 23716 6996
rect 25044 6944 25096 6996
rect 25596 6944 25648 6996
rect 23572 6876 23624 6928
rect 23204 6808 23256 6860
rect 18236 6740 18288 6792
rect 18696 6740 18748 6792
rect 21824 6672 21876 6724
rect 16580 6604 16632 6656
rect 18236 6604 18288 6656
rect 18788 6647 18840 6656
rect 18788 6613 18797 6647
rect 18797 6613 18831 6647
rect 18831 6613 18840 6647
rect 18788 6604 18840 6613
rect 22192 6740 22244 6792
rect 24952 6851 25004 6860
rect 24952 6817 24961 6851
rect 24961 6817 24995 6851
rect 24995 6817 25004 6851
rect 24952 6808 25004 6817
rect 23480 6740 23532 6792
rect 23756 6783 23808 6792
rect 23756 6749 23765 6783
rect 23765 6749 23799 6783
rect 23799 6749 23808 6783
rect 23756 6740 23808 6749
rect 22376 6672 22428 6724
rect 25688 6783 25740 6792
rect 25688 6749 25697 6783
rect 25697 6749 25731 6783
rect 25731 6749 25740 6783
rect 25688 6740 25740 6749
rect 22652 6647 22704 6656
rect 22652 6613 22661 6647
rect 22661 6613 22695 6647
rect 22695 6613 22704 6647
rect 22652 6604 22704 6613
rect 23296 6604 23348 6656
rect 25044 6604 25096 6656
rect 25136 6647 25188 6656
rect 25136 6613 25145 6647
rect 25145 6613 25179 6647
rect 25179 6613 25188 6647
rect 25136 6604 25188 6613
rect 25504 6604 25556 6656
rect 5083 6502 5135 6554
rect 5147 6502 5199 6554
rect 5211 6502 5263 6554
rect 5275 6502 5327 6554
rect 5339 6502 5391 6554
rect 12029 6502 12081 6554
rect 12093 6502 12145 6554
rect 12157 6502 12209 6554
rect 12221 6502 12273 6554
rect 12285 6502 12337 6554
rect 18975 6502 19027 6554
rect 19039 6502 19091 6554
rect 19103 6502 19155 6554
rect 19167 6502 19219 6554
rect 19231 6502 19283 6554
rect 25921 6502 25973 6554
rect 25985 6502 26037 6554
rect 26049 6502 26101 6554
rect 26113 6502 26165 6554
rect 26177 6502 26229 6554
rect 18236 6332 18288 6384
rect 19708 6332 19760 6384
rect 22192 6400 22244 6452
rect 22652 6443 22704 6452
rect 22652 6409 22661 6443
rect 22661 6409 22695 6443
rect 22695 6409 22704 6443
rect 22652 6400 22704 6409
rect 23204 6443 23256 6452
rect 23204 6409 23213 6443
rect 23213 6409 23247 6443
rect 23247 6409 23256 6443
rect 23204 6400 23256 6409
rect 23572 6400 23624 6452
rect 23756 6400 23808 6452
rect 22836 6375 22888 6384
rect 20536 6307 20588 6316
rect 20536 6273 20545 6307
rect 20545 6273 20579 6307
rect 20579 6273 20588 6307
rect 20536 6264 20588 6273
rect 20720 6264 20772 6316
rect 21180 6307 21232 6316
rect 21180 6273 21189 6307
rect 21189 6273 21223 6307
rect 21223 6273 21232 6307
rect 21180 6264 21232 6273
rect 22192 6264 22244 6316
rect 22836 6341 22845 6375
rect 22845 6341 22879 6375
rect 22879 6341 22888 6375
rect 22836 6332 22888 6341
rect 24768 6332 24820 6384
rect 24952 6332 25004 6384
rect 23020 6307 23072 6316
rect 23020 6273 23029 6307
rect 23029 6273 23063 6307
rect 23063 6273 23072 6307
rect 23020 6264 23072 6273
rect 23296 6264 23348 6316
rect 16580 6196 16632 6248
rect 17408 6196 17460 6248
rect 19340 6196 19392 6248
rect 22376 6128 22428 6180
rect 23480 6196 23532 6248
rect 23848 6264 23900 6316
rect 24032 6307 24084 6316
rect 24032 6273 24041 6307
rect 24041 6273 24075 6307
rect 24075 6273 24084 6307
rect 24032 6264 24084 6273
rect 28264 6307 28316 6316
rect 28264 6273 28273 6307
rect 28273 6273 28307 6307
rect 28307 6273 28316 6307
rect 28264 6264 28316 6273
rect 24216 6239 24268 6248
rect 24216 6205 24225 6239
rect 24225 6205 24259 6239
rect 24259 6205 24268 6239
rect 24216 6196 24268 6205
rect 24492 6239 24544 6248
rect 24492 6205 24501 6239
rect 24501 6205 24535 6239
rect 24535 6205 24544 6239
rect 24492 6196 24544 6205
rect 24584 6196 24636 6248
rect 25504 6196 25556 6248
rect 28540 6239 28592 6248
rect 28540 6205 28549 6239
rect 28549 6205 28583 6239
rect 28583 6205 28592 6239
rect 28540 6196 28592 6205
rect 19800 6060 19852 6112
rect 20168 6060 20220 6112
rect 22560 6060 22612 6112
rect 25044 6060 25096 6112
rect 4423 5958 4475 6010
rect 4487 5958 4539 6010
rect 4551 5958 4603 6010
rect 4615 5958 4667 6010
rect 4679 5958 4731 6010
rect 11369 5958 11421 6010
rect 11433 5958 11485 6010
rect 11497 5958 11549 6010
rect 11561 5958 11613 6010
rect 11625 5958 11677 6010
rect 18315 5958 18367 6010
rect 18379 5958 18431 6010
rect 18443 5958 18495 6010
rect 18507 5958 18559 6010
rect 18571 5958 18623 6010
rect 25261 5958 25313 6010
rect 25325 5958 25377 6010
rect 25389 5958 25441 6010
rect 25453 5958 25505 6010
rect 25517 5958 25569 6010
rect 20536 5856 20588 5908
rect 22744 5856 22796 5908
rect 24492 5856 24544 5908
rect 24584 5856 24636 5908
rect 25044 5856 25096 5908
rect 25136 5856 25188 5908
rect 19340 5788 19392 5840
rect 19800 5763 19852 5772
rect 19800 5729 19809 5763
rect 19809 5729 19843 5763
rect 19843 5729 19852 5763
rect 19800 5720 19852 5729
rect 17868 5652 17920 5704
rect 20076 5652 20128 5704
rect 20168 5695 20220 5704
rect 20168 5661 20177 5695
rect 20177 5661 20211 5695
rect 20211 5661 20220 5695
rect 20168 5652 20220 5661
rect 21732 5652 21784 5704
rect 23020 5720 23072 5772
rect 23940 5763 23992 5772
rect 23940 5729 23949 5763
rect 23949 5729 23983 5763
rect 23983 5729 23992 5763
rect 23940 5720 23992 5729
rect 22376 5695 22428 5704
rect 22376 5661 22385 5695
rect 22385 5661 22419 5695
rect 22419 5661 22428 5695
rect 22376 5652 22428 5661
rect 23664 5695 23716 5704
rect 23664 5661 23673 5695
rect 23673 5661 23707 5695
rect 23707 5661 23716 5695
rect 23664 5652 23716 5661
rect 23756 5695 23808 5704
rect 23756 5661 23765 5695
rect 23765 5661 23799 5695
rect 23799 5661 23808 5695
rect 23756 5652 23808 5661
rect 23848 5695 23900 5704
rect 23848 5661 23857 5695
rect 23857 5661 23891 5695
rect 23891 5661 23900 5695
rect 24768 5720 24820 5772
rect 23848 5652 23900 5661
rect 25688 5788 25740 5840
rect 16580 5516 16632 5568
rect 17960 5516 18012 5568
rect 19800 5516 19852 5568
rect 22100 5584 22152 5636
rect 22192 5584 22244 5636
rect 22284 5627 22336 5636
rect 22284 5593 22293 5627
rect 22293 5593 22327 5627
rect 22327 5593 22336 5627
rect 22284 5584 22336 5593
rect 22468 5627 22520 5636
rect 22468 5593 22503 5627
rect 22503 5593 22520 5627
rect 22468 5584 22520 5593
rect 24308 5584 24360 5636
rect 25596 5695 25648 5704
rect 25596 5661 25605 5695
rect 25605 5661 25639 5695
rect 25639 5661 25648 5695
rect 25596 5652 25648 5661
rect 5083 5414 5135 5466
rect 5147 5414 5199 5466
rect 5211 5414 5263 5466
rect 5275 5414 5327 5466
rect 5339 5414 5391 5466
rect 12029 5414 12081 5466
rect 12093 5414 12145 5466
rect 12157 5414 12209 5466
rect 12221 5414 12273 5466
rect 12285 5414 12337 5466
rect 18975 5414 19027 5466
rect 19039 5414 19091 5466
rect 19103 5414 19155 5466
rect 19167 5414 19219 5466
rect 19231 5414 19283 5466
rect 25921 5414 25973 5466
rect 25985 5414 26037 5466
rect 26049 5414 26101 5466
rect 26113 5414 26165 5466
rect 26177 5414 26229 5466
rect 18788 5244 18840 5296
rect 21916 5312 21968 5364
rect 22100 5312 22152 5364
rect 22192 5312 22244 5364
rect 22928 5355 22980 5364
rect 22928 5321 22937 5355
rect 22937 5321 22971 5355
rect 22971 5321 22980 5355
rect 22928 5312 22980 5321
rect 23204 5312 23256 5364
rect 16580 5108 16632 5160
rect 18236 5176 18288 5228
rect 19432 5176 19484 5228
rect 19892 5176 19944 5228
rect 20260 5176 20312 5228
rect 18328 5108 18380 5160
rect 20996 5176 21048 5228
rect 21640 5176 21692 5228
rect 18972 5040 19024 5092
rect 18052 4972 18104 5024
rect 19340 5015 19392 5024
rect 19340 4981 19349 5015
rect 19349 4981 19383 5015
rect 19383 4981 19392 5015
rect 19340 4972 19392 4981
rect 19708 4972 19760 5024
rect 20352 5015 20404 5024
rect 20352 4981 20361 5015
rect 20361 4981 20395 5015
rect 20395 4981 20404 5015
rect 20352 4972 20404 4981
rect 22284 5244 22336 5296
rect 22468 5040 22520 5092
rect 22284 4972 22336 5024
rect 22928 5176 22980 5228
rect 23756 5312 23808 5364
rect 23756 5219 23808 5228
rect 23756 5185 23765 5219
rect 23765 5185 23799 5219
rect 23799 5185 23808 5219
rect 23756 5176 23808 5185
rect 23940 5176 23992 5228
rect 24308 5219 24360 5228
rect 24308 5185 24317 5219
rect 24317 5185 24351 5219
rect 24351 5185 24360 5219
rect 24308 5176 24360 5185
rect 23020 5040 23072 5092
rect 24860 5176 24912 5228
rect 25596 5176 25648 5228
rect 25688 5176 25740 5228
rect 23756 4972 23808 5024
rect 24676 5015 24728 5024
rect 24676 4981 24685 5015
rect 24685 4981 24719 5015
rect 24719 4981 24728 5015
rect 24676 4972 24728 4981
rect 26148 4972 26200 5024
rect 4423 4870 4475 4922
rect 4487 4870 4539 4922
rect 4551 4870 4603 4922
rect 4615 4870 4667 4922
rect 4679 4870 4731 4922
rect 11369 4870 11421 4922
rect 11433 4870 11485 4922
rect 11497 4870 11549 4922
rect 11561 4870 11613 4922
rect 11625 4870 11677 4922
rect 18315 4870 18367 4922
rect 18379 4870 18431 4922
rect 18443 4870 18495 4922
rect 18507 4870 18559 4922
rect 18571 4870 18623 4922
rect 25261 4870 25313 4922
rect 25325 4870 25377 4922
rect 25389 4870 25441 4922
rect 25453 4870 25505 4922
rect 25517 4870 25569 4922
rect 17408 4768 17460 4820
rect 18236 4768 18288 4820
rect 19340 4768 19392 4820
rect 20996 4811 21048 4820
rect 20996 4777 21005 4811
rect 21005 4777 21039 4811
rect 21039 4777 21048 4811
rect 20996 4768 21048 4777
rect 22284 4768 22336 4820
rect 23296 4768 23348 4820
rect 24032 4768 24084 4820
rect 26148 4811 26200 4820
rect 26148 4777 26157 4811
rect 26157 4777 26191 4811
rect 26191 4777 26200 4811
rect 26148 4768 26200 4777
rect 16580 4632 16632 4684
rect 18880 4700 18932 4752
rect 17960 4607 18012 4616
rect 17960 4573 17969 4607
rect 17969 4573 18003 4607
rect 18003 4573 18012 4607
rect 17960 4564 18012 4573
rect 18788 4607 18840 4616
rect 18788 4573 18797 4607
rect 18797 4573 18831 4607
rect 18831 4573 18840 4607
rect 18788 4564 18840 4573
rect 18972 4564 19024 4616
rect 16120 4539 16172 4548
rect 16120 4505 16129 4539
rect 16129 4505 16163 4539
rect 16163 4505 16172 4539
rect 16120 4496 16172 4505
rect 17960 4428 18012 4480
rect 21272 4607 21324 4616
rect 21272 4573 21281 4607
rect 21281 4573 21315 4607
rect 21315 4573 21324 4607
rect 21272 4564 21324 4573
rect 21456 4607 21508 4616
rect 21456 4573 21465 4607
rect 21465 4573 21499 4607
rect 21499 4573 21508 4607
rect 21456 4564 21508 4573
rect 19524 4539 19576 4548
rect 19524 4505 19533 4539
rect 19533 4505 19567 4539
rect 19567 4505 19576 4539
rect 19524 4496 19576 4505
rect 19616 4496 19668 4548
rect 19800 4428 19852 4480
rect 21548 4428 21600 4480
rect 22744 4607 22796 4616
rect 22744 4573 22753 4607
rect 22753 4573 22787 4607
rect 22787 4573 22796 4607
rect 22744 4564 22796 4573
rect 22836 4539 22888 4548
rect 22836 4505 22845 4539
rect 22845 4505 22879 4539
rect 22879 4505 22888 4539
rect 22836 4496 22888 4505
rect 24216 4632 24268 4684
rect 24676 4675 24728 4684
rect 24676 4641 24685 4675
rect 24685 4641 24719 4675
rect 24719 4641 24728 4675
rect 24676 4632 24728 4641
rect 23112 4496 23164 4548
rect 24952 4496 25004 4548
rect 25136 4496 25188 4548
rect 21916 4471 21968 4480
rect 21916 4437 21925 4471
rect 21925 4437 21959 4471
rect 21959 4437 21968 4471
rect 21916 4428 21968 4437
rect 22652 4471 22704 4480
rect 22652 4437 22661 4471
rect 22661 4437 22695 4471
rect 22695 4437 22704 4471
rect 22652 4428 22704 4437
rect 22928 4471 22980 4480
rect 22928 4437 22937 4471
rect 22937 4437 22971 4471
rect 22971 4437 22980 4471
rect 22928 4428 22980 4437
rect 23296 4428 23348 4480
rect 23480 4428 23532 4480
rect 5083 4326 5135 4378
rect 5147 4326 5199 4378
rect 5211 4326 5263 4378
rect 5275 4326 5327 4378
rect 5339 4326 5391 4378
rect 12029 4326 12081 4378
rect 12093 4326 12145 4378
rect 12157 4326 12209 4378
rect 12221 4326 12273 4378
rect 12285 4326 12337 4378
rect 18975 4326 19027 4378
rect 19039 4326 19091 4378
rect 19103 4326 19155 4378
rect 19167 4326 19219 4378
rect 19231 4326 19283 4378
rect 25921 4326 25973 4378
rect 25985 4326 26037 4378
rect 26049 4326 26101 4378
rect 26113 4326 26165 4378
rect 26177 4326 26229 4378
rect 16120 4224 16172 4276
rect 19524 4224 19576 4276
rect 20352 4224 20404 4276
rect 21548 4267 21600 4276
rect 21548 4233 21557 4267
rect 21557 4233 21591 4267
rect 21591 4233 21600 4267
rect 21548 4224 21600 4233
rect 21916 4224 21968 4276
rect 17132 4088 17184 4140
rect 18972 4131 19024 4140
rect 18972 4097 18981 4131
rect 18981 4097 19015 4131
rect 19015 4097 19024 4131
rect 18972 4088 19024 4097
rect 19340 4131 19392 4140
rect 19340 4097 19349 4131
rect 19349 4097 19383 4131
rect 19383 4097 19392 4131
rect 19340 4088 19392 4097
rect 19432 4088 19484 4140
rect 18052 4020 18104 4072
rect 18696 4020 18748 4072
rect 17408 3884 17460 3936
rect 21732 4156 21784 4208
rect 22468 4224 22520 4276
rect 23020 4224 23072 4276
rect 23572 4224 23624 4276
rect 24032 4224 24084 4276
rect 24952 4267 25004 4276
rect 24952 4233 24961 4267
rect 24961 4233 24995 4267
rect 24995 4233 25004 4267
rect 24952 4224 25004 4233
rect 22192 4199 22244 4208
rect 22192 4165 22201 4199
rect 22201 4165 22235 4199
rect 22235 4165 22244 4199
rect 22192 4156 22244 4165
rect 19800 4063 19852 4072
rect 19800 4029 19809 4063
rect 19809 4029 19843 4063
rect 19843 4029 19852 4063
rect 19800 4020 19852 4029
rect 22652 4088 22704 4140
rect 22836 4131 22888 4140
rect 22836 4097 22845 4131
rect 22845 4097 22879 4131
rect 22879 4097 22888 4131
rect 22836 4088 22888 4097
rect 23020 4088 23072 4140
rect 23112 4088 23164 4140
rect 22928 3952 22980 4004
rect 23572 4088 23624 4140
rect 24768 4020 24820 4072
rect 26148 4020 26200 4072
rect 19708 3884 19760 3936
rect 20260 3884 20312 3936
rect 23388 3927 23440 3936
rect 23388 3893 23397 3927
rect 23397 3893 23431 3927
rect 23431 3893 23440 3927
rect 23388 3884 23440 3893
rect 23664 3927 23716 3936
rect 23664 3893 23673 3927
rect 23673 3893 23707 3927
rect 23707 3893 23716 3927
rect 23664 3884 23716 3893
rect 23756 3927 23808 3936
rect 23756 3893 23765 3927
rect 23765 3893 23799 3927
rect 23799 3893 23808 3927
rect 23756 3884 23808 3893
rect 4423 3782 4475 3834
rect 4487 3782 4539 3834
rect 4551 3782 4603 3834
rect 4615 3782 4667 3834
rect 4679 3782 4731 3834
rect 11369 3782 11421 3834
rect 11433 3782 11485 3834
rect 11497 3782 11549 3834
rect 11561 3782 11613 3834
rect 11625 3782 11677 3834
rect 18315 3782 18367 3834
rect 18379 3782 18431 3834
rect 18443 3782 18495 3834
rect 18507 3782 18559 3834
rect 18571 3782 18623 3834
rect 25261 3782 25313 3834
rect 25325 3782 25377 3834
rect 25389 3782 25441 3834
rect 25453 3782 25505 3834
rect 25517 3782 25569 3834
rect 19432 3680 19484 3732
rect 16580 3587 16632 3596
rect 16580 3553 16589 3587
rect 16589 3553 16623 3587
rect 16623 3553 16632 3587
rect 16580 3544 16632 3553
rect 19616 3544 19668 3596
rect 19892 3587 19944 3596
rect 19892 3553 19901 3587
rect 19901 3553 19935 3587
rect 19935 3553 19944 3587
rect 19892 3544 19944 3553
rect 21456 3680 21508 3732
rect 22192 3680 22244 3732
rect 22744 3680 22796 3732
rect 23020 3680 23072 3732
rect 23388 3680 23440 3732
rect 26148 3723 26200 3732
rect 26148 3689 26157 3723
rect 26157 3689 26191 3723
rect 26191 3689 26200 3723
rect 26148 3680 26200 3689
rect 17868 3476 17920 3528
rect 17960 3476 18012 3528
rect 18604 3476 18656 3528
rect 20260 3519 20312 3528
rect 20260 3485 20269 3519
rect 20269 3485 20303 3519
rect 20303 3485 20312 3519
rect 20260 3476 20312 3485
rect 20812 3519 20864 3528
rect 20812 3485 20821 3519
rect 20821 3485 20855 3519
rect 20855 3485 20864 3519
rect 20812 3476 20864 3485
rect 16856 3451 16908 3460
rect 16856 3417 16865 3451
rect 16865 3417 16899 3451
rect 16899 3417 16908 3451
rect 16856 3408 16908 3417
rect 20904 3408 20956 3460
rect 18880 3340 18932 3392
rect 19340 3340 19392 3392
rect 20720 3383 20772 3392
rect 20720 3349 20729 3383
rect 20729 3349 20763 3383
rect 20763 3349 20772 3383
rect 20720 3340 20772 3349
rect 21824 3340 21876 3392
rect 24216 3544 24268 3596
rect 22560 3408 22612 3460
rect 22652 3383 22704 3392
rect 22652 3349 22661 3383
rect 22661 3349 22695 3383
rect 22695 3349 22704 3383
rect 22652 3340 22704 3349
rect 23112 3408 23164 3460
rect 23296 3519 23348 3528
rect 23296 3485 23305 3519
rect 23305 3485 23339 3519
rect 23339 3485 23348 3519
rect 23296 3476 23348 3485
rect 23480 3476 23532 3528
rect 23756 3476 23808 3528
rect 25136 3408 25188 3460
rect 23296 3340 23348 3392
rect 5083 3238 5135 3290
rect 5147 3238 5199 3290
rect 5211 3238 5263 3290
rect 5275 3238 5327 3290
rect 5339 3238 5391 3290
rect 12029 3238 12081 3290
rect 12093 3238 12145 3290
rect 12157 3238 12209 3290
rect 12221 3238 12273 3290
rect 12285 3238 12337 3290
rect 18975 3238 19027 3290
rect 19039 3238 19091 3290
rect 19103 3238 19155 3290
rect 19167 3238 19219 3290
rect 19231 3238 19283 3290
rect 25921 3238 25973 3290
rect 25985 3238 26037 3290
rect 26049 3238 26101 3290
rect 26113 3238 26165 3290
rect 26177 3238 26229 3290
rect 16856 3136 16908 3188
rect 17408 3136 17460 3188
rect 19524 3136 19576 3188
rect 19616 3179 19668 3188
rect 19616 3145 19625 3179
rect 19625 3145 19659 3179
rect 19659 3145 19668 3179
rect 19616 3136 19668 3145
rect 18604 3068 18656 3120
rect 17868 3043 17920 3052
rect 17868 3009 17877 3043
rect 17877 3009 17911 3043
rect 17911 3009 17920 3043
rect 17868 3000 17920 3009
rect 19800 3136 19852 3188
rect 21732 3068 21784 3120
rect 19984 2975 20036 2984
rect 19984 2941 19993 2975
rect 19993 2941 20027 2975
rect 20027 2941 20036 2975
rect 19984 2932 20036 2941
rect 21180 2932 21232 2984
rect 21456 2907 21508 2916
rect 21456 2873 21465 2907
rect 21465 2873 21499 2907
rect 21499 2873 21508 2907
rect 21456 2864 21508 2873
rect 21824 3043 21876 3052
rect 21824 3009 21833 3043
rect 21833 3009 21867 3043
rect 21867 3009 21876 3043
rect 21824 3000 21876 3009
rect 22100 2975 22152 2984
rect 22100 2941 22109 2975
rect 22109 2941 22143 2975
rect 22143 2941 22152 2975
rect 22100 2932 22152 2941
rect 25136 3000 25188 3052
rect 23480 2932 23532 2984
rect 23664 2839 23716 2848
rect 23664 2805 23673 2839
rect 23673 2805 23707 2839
rect 23707 2805 23716 2839
rect 23664 2796 23716 2805
rect 4423 2694 4475 2746
rect 4487 2694 4539 2746
rect 4551 2694 4603 2746
rect 4615 2694 4667 2746
rect 4679 2694 4731 2746
rect 11369 2694 11421 2746
rect 11433 2694 11485 2746
rect 11497 2694 11549 2746
rect 11561 2694 11613 2746
rect 11625 2694 11677 2746
rect 18315 2694 18367 2746
rect 18379 2694 18431 2746
rect 18443 2694 18495 2746
rect 18507 2694 18559 2746
rect 18571 2694 18623 2746
rect 25261 2694 25313 2746
rect 25325 2694 25377 2746
rect 25389 2694 25441 2746
rect 25453 2694 25505 2746
rect 25517 2694 25569 2746
rect 18144 2635 18196 2644
rect 18144 2601 18153 2635
rect 18153 2601 18187 2635
rect 18187 2601 18196 2635
rect 18144 2592 18196 2601
rect 19984 2592 20036 2644
rect 21180 2635 21232 2644
rect 21180 2601 21189 2635
rect 21189 2601 21223 2635
rect 21223 2601 21232 2635
rect 21180 2592 21232 2601
rect 21272 2592 21324 2644
rect 22100 2592 22152 2644
rect 23296 2592 23348 2644
rect 13544 2456 13596 2508
rect 19340 2499 19392 2508
rect 19340 2465 19349 2499
rect 19349 2465 19383 2499
rect 19383 2465 19392 2499
rect 19340 2456 19392 2465
rect 22652 2499 22704 2508
rect 22652 2465 22661 2499
rect 22661 2465 22695 2499
rect 22695 2465 22704 2499
rect 22652 2456 22704 2465
rect 20 2388 72 2440
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 18052 2388 18104 2440
rect 19616 2388 19668 2440
rect 20720 2388 20772 2440
rect 20904 2388 20956 2440
rect 23664 2456 23716 2508
rect 17132 2320 17184 2372
rect 23112 2388 23164 2440
rect 23388 2388 23440 2440
rect 27068 2388 27120 2440
rect 18788 2252 18840 2304
rect 5083 2150 5135 2202
rect 5147 2150 5199 2202
rect 5211 2150 5263 2202
rect 5275 2150 5327 2202
rect 5339 2150 5391 2202
rect 12029 2150 12081 2202
rect 12093 2150 12145 2202
rect 12157 2150 12209 2202
rect 12221 2150 12273 2202
rect 12285 2150 12337 2202
rect 18975 2150 19027 2202
rect 19039 2150 19091 2202
rect 19103 2150 19155 2202
rect 19167 2150 19219 2202
rect 19231 2150 19283 2202
rect 25921 2150 25973 2202
rect 25985 2150 26037 2202
rect 26049 2150 26101 2202
rect 26113 2150 26165 2202
rect 26177 2150 26229 2202
<< metal2 >>
rect 7102 29322 7158 30000
rect 7102 29294 7236 29322
rect 7102 29200 7158 29294
rect 4423 27772 4731 27781
rect 4423 27770 4429 27772
rect 4485 27770 4509 27772
rect 4565 27770 4589 27772
rect 4645 27770 4669 27772
rect 4725 27770 4731 27772
rect 4485 27718 4487 27770
rect 4667 27718 4669 27770
rect 4423 27716 4429 27718
rect 4485 27716 4509 27718
rect 4565 27716 4589 27718
rect 4645 27716 4669 27718
rect 4725 27716 4731 27718
rect 1490 27704 1546 27713
rect 4423 27707 4731 27716
rect 1490 27639 1546 27648
rect 1504 27606 1532 27639
rect 7208 27606 7236 29294
rect 16118 29200 16174 30000
rect 25134 29200 25190 30000
rect 11369 27772 11677 27781
rect 11369 27770 11375 27772
rect 11431 27770 11455 27772
rect 11511 27770 11535 27772
rect 11591 27770 11615 27772
rect 11671 27770 11677 27772
rect 11431 27718 11433 27770
rect 11613 27718 11615 27770
rect 11369 27716 11375 27718
rect 11431 27716 11455 27718
rect 11511 27716 11535 27718
rect 11591 27716 11615 27718
rect 11671 27716 11677 27718
rect 11369 27707 11677 27716
rect 16132 27606 16160 29200
rect 18315 27772 18623 27781
rect 18315 27770 18321 27772
rect 18377 27770 18401 27772
rect 18457 27770 18481 27772
rect 18537 27770 18561 27772
rect 18617 27770 18623 27772
rect 18377 27718 18379 27770
rect 18559 27718 18561 27770
rect 18315 27716 18321 27718
rect 18377 27716 18401 27718
rect 18457 27716 18481 27718
rect 18537 27716 18561 27718
rect 18617 27716 18623 27718
rect 18315 27707 18623 27716
rect 1492 27600 1544 27606
rect 1492 27542 1544 27548
rect 7196 27600 7248 27606
rect 7196 27542 7248 27548
rect 16120 27600 16172 27606
rect 16120 27542 16172 27548
rect 21640 27600 21692 27606
rect 21640 27542 21692 27548
rect 17592 27464 17644 27470
rect 17592 27406 17644 27412
rect 15844 27328 15896 27334
rect 15844 27270 15896 27276
rect 5083 27228 5391 27237
rect 5083 27226 5089 27228
rect 5145 27226 5169 27228
rect 5225 27226 5249 27228
rect 5305 27226 5329 27228
rect 5385 27226 5391 27228
rect 5145 27174 5147 27226
rect 5327 27174 5329 27226
rect 5083 27172 5089 27174
rect 5145 27172 5169 27174
rect 5225 27172 5249 27174
rect 5305 27172 5329 27174
rect 5385 27172 5391 27174
rect 5083 27163 5391 27172
rect 12029 27228 12337 27237
rect 12029 27226 12035 27228
rect 12091 27226 12115 27228
rect 12171 27226 12195 27228
rect 12251 27226 12275 27228
rect 12331 27226 12337 27228
rect 12091 27174 12093 27226
rect 12273 27174 12275 27226
rect 12029 27172 12035 27174
rect 12091 27172 12115 27174
rect 12171 27172 12195 27174
rect 12251 27172 12275 27174
rect 12331 27172 12337 27174
rect 12029 27163 12337 27172
rect 4423 26684 4731 26693
rect 4423 26682 4429 26684
rect 4485 26682 4509 26684
rect 4565 26682 4589 26684
rect 4645 26682 4669 26684
rect 4725 26682 4731 26684
rect 4485 26630 4487 26682
rect 4667 26630 4669 26682
rect 4423 26628 4429 26630
rect 4485 26628 4509 26630
rect 4565 26628 4589 26630
rect 4645 26628 4669 26630
rect 4725 26628 4731 26630
rect 4423 26619 4731 26628
rect 11369 26684 11677 26693
rect 11369 26682 11375 26684
rect 11431 26682 11455 26684
rect 11511 26682 11535 26684
rect 11591 26682 11615 26684
rect 11671 26682 11677 26684
rect 11431 26630 11433 26682
rect 11613 26630 11615 26682
rect 11369 26628 11375 26630
rect 11431 26628 11455 26630
rect 11511 26628 11535 26630
rect 11591 26628 11615 26630
rect 11671 26628 11677 26630
rect 11369 26619 11677 26628
rect 5083 26140 5391 26149
rect 5083 26138 5089 26140
rect 5145 26138 5169 26140
rect 5225 26138 5249 26140
rect 5305 26138 5329 26140
rect 5385 26138 5391 26140
rect 5145 26086 5147 26138
rect 5327 26086 5329 26138
rect 5083 26084 5089 26086
rect 5145 26084 5169 26086
rect 5225 26084 5249 26086
rect 5305 26084 5329 26086
rect 5385 26084 5391 26086
rect 5083 26075 5391 26084
rect 12029 26140 12337 26149
rect 12029 26138 12035 26140
rect 12091 26138 12115 26140
rect 12171 26138 12195 26140
rect 12251 26138 12275 26140
rect 12331 26138 12337 26140
rect 12091 26086 12093 26138
rect 12273 26086 12275 26138
rect 12029 26084 12035 26086
rect 12091 26084 12115 26086
rect 12171 26084 12195 26086
rect 12251 26084 12275 26086
rect 12331 26084 12337 26086
rect 12029 26075 12337 26084
rect 4423 25596 4731 25605
rect 4423 25594 4429 25596
rect 4485 25594 4509 25596
rect 4565 25594 4589 25596
rect 4645 25594 4669 25596
rect 4725 25594 4731 25596
rect 4485 25542 4487 25594
rect 4667 25542 4669 25594
rect 4423 25540 4429 25542
rect 4485 25540 4509 25542
rect 4565 25540 4589 25542
rect 4645 25540 4669 25542
rect 4725 25540 4731 25542
rect 4423 25531 4731 25540
rect 11369 25596 11677 25605
rect 11369 25594 11375 25596
rect 11431 25594 11455 25596
rect 11511 25594 11535 25596
rect 11591 25594 11615 25596
rect 11671 25594 11677 25596
rect 11431 25542 11433 25594
rect 11613 25542 11615 25594
rect 11369 25540 11375 25542
rect 11431 25540 11455 25542
rect 11511 25540 11535 25542
rect 11591 25540 11615 25542
rect 11671 25540 11677 25542
rect 11369 25531 11677 25540
rect 5083 25052 5391 25061
rect 5083 25050 5089 25052
rect 5145 25050 5169 25052
rect 5225 25050 5249 25052
rect 5305 25050 5329 25052
rect 5385 25050 5391 25052
rect 5145 24998 5147 25050
rect 5327 24998 5329 25050
rect 5083 24996 5089 24998
rect 5145 24996 5169 24998
rect 5225 24996 5249 24998
rect 5305 24996 5329 24998
rect 5385 24996 5391 24998
rect 5083 24987 5391 24996
rect 12029 25052 12337 25061
rect 12029 25050 12035 25052
rect 12091 25050 12115 25052
rect 12171 25050 12195 25052
rect 12251 25050 12275 25052
rect 12331 25050 12337 25052
rect 12091 24998 12093 25050
rect 12273 24998 12275 25050
rect 12029 24996 12035 24998
rect 12091 24996 12115 24998
rect 12171 24996 12195 24998
rect 12251 24996 12275 24998
rect 12331 24996 12337 24998
rect 12029 24987 12337 24996
rect 4423 24508 4731 24517
rect 4423 24506 4429 24508
rect 4485 24506 4509 24508
rect 4565 24506 4589 24508
rect 4645 24506 4669 24508
rect 4725 24506 4731 24508
rect 4485 24454 4487 24506
rect 4667 24454 4669 24506
rect 4423 24452 4429 24454
rect 4485 24452 4509 24454
rect 4565 24452 4589 24454
rect 4645 24452 4669 24454
rect 4725 24452 4731 24454
rect 4423 24443 4731 24452
rect 11369 24508 11677 24517
rect 11369 24506 11375 24508
rect 11431 24506 11455 24508
rect 11511 24506 11535 24508
rect 11591 24506 11615 24508
rect 11671 24506 11677 24508
rect 11431 24454 11433 24506
rect 11613 24454 11615 24506
rect 11369 24452 11375 24454
rect 11431 24452 11455 24454
rect 11511 24452 11535 24454
rect 11591 24452 11615 24454
rect 11671 24452 11677 24454
rect 11369 24443 11677 24452
rect 5083 23964 5391 23973
rect 5083 23962 5089 23964
rect 5145 23962 5169 23964
rect 5225 23962 5249 23964
rect 5305 23962 5329 23964
rect 5385 23962 5391 23964
rect 5145 23910 5147 23962
rect 5327 23910 5329 23962
rect 5083 23908 5089 23910
rect 5145 23908 5169 23910
rect 5225 23908 5249 23910
rect 5305 23908 5329 23910
rect 5385 23908 5391 23910
rect 5083 23899 5391 23908
rect 12029 23964 12337 23973
rect 12029 23962 12035 23964
rect 12091 23962 12115 23964
rect 12171 23962 12195 23964
rect 12251 23962 12275 23964
rect 12331 23962 12337 23964
rect 12091 23910 12093 23962
rect 12273 23910 12275 23962
rect 12029 23908 12035 23910
rect 12091 23908 12115 23910
rect 12171 23908 12195 23910
rect 12251 23908 12275 23910
rect 12331 23908 12337 23910
rect 12029 23899 12337 23908
rect 4423 23420 4731 23429
rect 4423 23418 4429 23420
rect 4485 23418 4509 23420
rect 4565 23418 4589 23420
rect 4645 23418 4669 23420
rect 4725 23418 4731 23420
rect 4485 23366 4487 23418
rect 4667 23366 4669 23418
rect 4423 23364 4429 23366
rect 4485 23364 4509 23366
rect 4565 23364 4589 23366
rect 4645 23364 4669 23366
rect 4725 23364 4731 23366
rect 4423 23355 4731 23364
rect 11369 23420 11677 23429
rect 11369 23418 11375 23420
rect 11431 23418 11455 23420
rect 11511 23418 11535 23420
rect 11591 23418 11615 23420
rect 11671 23418 11677 23420
rect 11431 23366 11433 23418
rect 11613 23366 11615 23418
rect 11369 23364 11375 23366
rect 11431 23364 11455 23366
rect 11511 23364 11535 23366
rect 11591 23364 11615 23366
rect 11671 23364 11677 23366
rect 11369 23355 11677 23364
rect 5083 22876 5391 22885
rect 5083 22874 5089 22876
rect 5145 22874 5169 22876
rect 5225 22874 5249 22876
rect 5305 22874 5329 22876
rect 5385 22874 5391 22876
rect 5145 22822 5147 22874
rect 5327 22822 5329 22874
rect 5083 22820 5089 22822
rect 5145 22820 5169 22822
rect 5225 22820 5249 22822
rect 5305 22820 5329 22822
rect 5385 22820 5391 22822
rect 5083 22811 5391 22820
rect 12029 22876 12337 22885
rect 12029 22874 12035 22876
rect 12091 22874 12115 22876
rect 12171 22874 12195 22876
rect 12251 22874 12275 22876
rect 12331 22874 12337 22876
rect 12091 22822 12093 22874
rect 12273 22822 12275 22874
rect 12029 22820 12035 22822
rect 12091 22820 12115 22822
rect 12171 22820 12195 22822
rect 12251 22820 12275 22822
rect 12331 22820 12337 22822
rect 12029 22811 12337 22820
rect 4423 22332 4731 22341
rect 4423 22330 4429 22332
rect 4485 22330 4509 22332
rect 4565 22330 4589 22332
rect 4645 22330 4669 22332
rect 4725 22330 4731 22332
rect 4485 22278 4487 22330
rect 4667 22278 4669 22330
rect 4423 22276 4429 22278
rect 4485 22276 4509 22278
rect 4565 22276 4589 22278
rect 4645 22276 4669 22278
rect 4725 22276 4731 22278
rect 4423 22267 4731 22276
rect 11369 22332 11677 22341
rect 11369 22330 11375 22332
rect 11431 22330 11455 22332
rect 11511 22330 11535 22332
rect 11591 22330 11615 22332
rect 11671 22330 11677 22332
rect 11431 22278 11433 22330
rect 11613 22278 11615 22330
rect 11369 22276 11375 22278
rect 11431 22276 11455 22278
rect 11511 22276 11535 22278
rect 11591 22276 11615 22278
rect 11671 22276 11677 22278
rect 11369 22267 11677 22276
rect 5083 21788 5391 21797
rect 5083 21786 5089 21788
rect 5145 21786 5169 21788
rect 5225 21786 5249 21788
rect 5305 21786 5329 21788
rect 5385 21786 5391 21788
rect 5145 21734 5147 21786
rect 5327 21734 5329 21786
rect 5083 21732 5089 21734
rect 5145 21732 5169 21734
rect 5225 21732 5249 21734
rect 5305 21732 5329 21734
rect 5385 21732 5391 21734
rect 5083 21723 5391 21732
rect 12029 21788 12337 21797
rect 12029 21786 12035 21788
rect 12091 21786 12115 21788
rect 12171 21786 12195 21788
rect 12251 21786 12275 21788
rect 12331 21786 12337 21788
rect 12091 21734 12093 21786
rect 12273 21734 12275 21786
rect 12029 21732 12035 21734
rect 12091 21732 12115 21734
rect 12171 21732 12195 21734
rect 12251 21732 12275 21734
rect 12331 21732 12337 21734
rect 12029 21723 12337 21732
rect 4423 21244 4731 21253
rect 4423 21242 4429 21244
rect 4485 21242 4509 21244
rect 4565 21242 4589 21244
rect 4645 21242 4669 21244
rect 4725 21242 4731 21244
rect 4485 21190 4487 21242
rect 4667 21190 4669 21242
rect 4423 21188 4429 21190
rect 4485 21188 4509 21190
rect 4565 21188 4589 21190
rect 4645 21188 4669 21190
rect 4725 21188 4731 21190
rect 4423 21179 4731 21188
rect 11369 21244 11677 21253
rect 11369 21242 11375 21244
rect 11431 21242 11455 21244
rect 11511 21242 11535 21244
rect 11591 21242 11615 21244
rect 11671 21242 11677 21244
rect 11431 21190 11433 21242
rect 11613 21190 11615 21242
rect 11369 21188 11375 21190
rect 11431 21188 11455 21190
rect 11511 21188 11535 21190
rect 11591 21188 11615 21190
rect 11671 21188 11677 21190
rect 11369 21179 11677 21188
rect 5083 20700 5391 20709
rect 5083 20698 5089 20700
rect 5145 20698 5169 20700
rect 5225 20698 5249 20700
rect 5305 20698 5329 20700
rect 5385 20698 5391 20700
rect 5145 20646 5147 20698
rect 5327 20646 5329 20698
rect 5083 20644 5089 20646
rect 5145 20644 5169 20646
rect 5225 20644 5249 20646
rect 5305 20644 5329 20646
rect 5385 20644 5391 20646
rect 5083 20635 5391 20644
rect 12029 20700 12337 20709
rect 12029 20698 12035 20700
rect 12091 20698 12115 20700
rect 12171 20698 12195 20700
rect 12251 20698 12275 20700
rect 12331 20698 12337 20700
rect 12091 20646 12093 20698
rect 12273 20646 12275 20698
rect 12029 20644 12035 20646
rect 12091 20644 12115 20646
rect 12171 20644 12195 20646
rect 12251 20644 12275 20646
rect 12331 20644 12337 20646
rect 12029 20635 12337 20644
rect 4423 20156 4731 20165
rect 4423 20154 4429 20156
rect 4485 20154 4509 20156
rect 4565 20154 4589 20156
rect 4645 20154 4669 20156
rect 4725 20154 4731 20156
rect 4485 20102 4487 20154
rect 4667 20102 4669 20154
rect 4423 20100 4429 20102
rect 4485 20100 4509 20102
rect 4565 20100 4589 20102
rect 4645 20100 4669 20102
rect 4725 20100 4731 20102
rect 4423 20091 4731 20100
rect 11369 20156 11677 20165
rect 11369 20154 11375 20156
rect 11431 20154 11455 20156
rect 11511 20154 11535 20156
rect 11591 20154 11615 20156
rect 11671 20154 11677 20156
rect 11431 20102 11433 20154
rect 11613 20102 11615 20154
rect 11369 20100 11375 20102
rect 11431 20100 11455 20102
rect 11511 20100 11535 20102
rect 11591 20100 11615 20102
rect 11671 20100 11677 20102
rect 11369 20091 11677 20100
rect 5083 19612 5391 19621
rect 5083 19610 5089 19612
rect 5145 19610 5169 19612
rect 5225 19610 5249 19612
rect 5305 19610 5329 19612
rect 5385 19610 5391 19612
rect 5145 19558 5147 19610
rect 5327 19558 5329 19610
rect 5083 19556 5089 19558
rect 5145 19556 5169 19558
rect 5225 19556 5249 19558
rect 5305 19556 5329 19558
rect 5385 19556 5391 19558
rect 5083 19547 5391 19556
rect 12029 19612 12337 19621
rect 12029 19610 12035 19612
rect 12091 19610 12115 19612
rect 12171 19610 12195 19612
rect 12251 19610 12275 19612
rect 12331 19610 12337 19612
rect 12091 19558 12093 19610
rect 12273 19558 12275 19610
rect 12029 19556 12035 19558
rect 12091 19556 12115 19558
rect 12171 19556 12195 19558
rect 12251 19556 12275 19558
rect 12331 19556 12337 19558
rect 12029 19547 12337 19556
rect 4423 19068 4731 19077
rect 4423 19066 4429 19068
rect 4485 19066 4509 19068
rect 4565 19066 4589 19068
rect 4645 19066 4669 19068
rect 4725 19066 4731 19068
rect 4485 19014 4487 19066
rect 4667 19014 4669 19066
rect 4423 19012 4429 19014
rect 4485 19012 4509 19014
rect 4565 19012 4589 19014
rect 4645 19012 4669 19014
rect 4725 19012 4731 19014
rect 4423 19003 4731 19012
rect 11369 19068 11677 19077
rect 11369 19066 11375 19068
rect 11431 19066 11455 19068
rect 11511 19066 11535 19068
rect 11591 19066 11615 19068
rect 11671 19066 11677 19068
rect 11431 19014 11433 19066
rect 11613 19014 11615 19066
rect 11369 19012 11375 19014
rect 11431 19012 11455 19014
rect 11511 19012 11535 19014
rect 11591 19012 11615 19014
rect 11671 19012 11677 19014
rect 11369 19003 11677 19012
rect 940 18760 992 18766
rect 940 18702 992 18708
rect 13452 18760 13504 18766
rect 13452 18702 13504 18708
rect 952 18465 980 18702
rect 5083 18524 5391 18533
rect 5083 18522 5089 18524
rect 5145 18522 5169 18524
rect 5225 18522 5249 18524
rect 5305 18522 5329 18524
rect 5385 18522 5391 18524
rect 5145 18470 5147 18522
rect 5327 18470 5329 18522
rect 5083 18468 5089 18470
rect 5145 18468 5169 18470
rect 5225 18468 5249 18470
rect 5305 18468 5329 18470
rect 5385 18468 5391 18470
rect 938 18456 994 18465
rect 5083 18459 5391 18468
rect 12029 18524 12337 18533
rect 12029 18522 12035 18524
rect 12091 18522 12115 18524
rect 12171 18522 12195 18524
rect 12251 18522 12275 18524
rect 12331 18522 12337 18524
rect 12091 18470 12093 18522
rect 12273 18470 12275 18522
rect 12029 18468 12035 18470
rect 12091 18468 12115 18470
rect 12171 18468 12195 18470
rect 12251 18468 12275 18470
rect 12331 18468 12337 18470
rect 12029 18459 12337 18468
rect 938 18391 994 18400
rect 4423 17980 4731 17989
rect 4423 17978 4429 17980
rect 4485 17978 4509 17980
rect 4565 17978 4589 17980
rect 4645 17978 4669 17980
rect 4725 17978 4731 17980
rect 4485 17926 4487 17978
rect 4667 17926 4669 17978
rect 4423 17924 4429 17926
rect 4485 17924 4509 17926
rect 4565 17924 4589 17926
rect 4645 17924 4669 17926
rect 4725 17924 4731 17926
rect 4423 17915 4731 17924
rect 11369 17980 11677 17989
rect 11369 17978 11375 17980
rect 11431 17978 11455 17980
rect 11511 17978 11535 17980
rect 11591 17978 11615 17980
rect 11671 17978 11677 17980
rect 11431 17926 11433 17978
rect 11613 17926 11615 17978
rect 11369 17924 11375 17926
rect 11431 17924 11455 17926
rect 11511 17924 11535 17926
rect 11591 17924 11615 17926
rect 11671 17924 11677 17926
rect 11369 17915 11677 17924
rect 5083 17436 5391 17445
rect 5083 17434 5089 17436
rect 5145 17434 5169 17436
rect 5225 17434 5249 17436
rect 5305 17434 5329 17436
rect 5385 17434 5391 17436
rect 5145 17382 5147 17434
rect 5327 17382 5329 17434
rect 5083 17380 5089 17382
rect 5145 17380 5169 17382
rect 5225 17380 5249 17382
rect 5305 17380 5329 17382
rect 5385 17380 5391 17382
rect 5083 17371 5391 17380
rect 12029 17436 12337 17445
rect 12029 17434 12035 17436
rect 12091 17434 12115 17436
rect 12171 17434 12195 17436
rect 12251 17434 12275 17436
rect 12331 17434 12337 17436
rect 12091 17382 12093 17434
rect 12273 17382 12275 17434
rect 12029 17380 12035 17382
rect 12091 17380 12115 17382
rect 12171 17380 12195 17382
rect 12251 17380 12275 17382
rect 12331 17380 12337 17382
rect 12029 17371 12337 17380
rect 4423 16892 4731 16901
rect 4423 16890 4429 16892
rect 4485 16890 4509 16892
rect 4565 16890 4589 16892
rect 4645 16890 4669 16892
rect 4725 16890 4731 16892
rect 4485 16838 4487 16890
rect 4667 16838 4669 16890
rect 4423 16836 4429 16838
rect 4485 16836 4509 16838
rect 4565 16836 4589 16838
rect 4645 16836 4669 16838
rect 4725 16836 4731 16838
rect 4423 16827 4731 16836
rect 11369 16892 11677 16901
rect 11369 16890 11375 16892
rect 11431 16890 11455 16892
rect 11511 16890 11535 16892
rect 11591 16890 11615 16892
rect 11671 16890 11677 16892
rect 11431 16838 11433 16890
rect 11613 16838 11615 16890
rect 11369 16836 11375 16838
rect 11431 16836 11455 16838
rect 11511 16836 11535 16838
rect 11591 16836 11615 16838
rect 11671 16836 11677 16838
rect 11369 16827 11677 16836
rect 5083 16348 5391 16357
rect 5083 16346 5089 16348
rect 5145 16346 5169 16348
rect 5225 16346 5249 16348
rect 5305 16346 5329 16348
rect 5385 16346 5391 16348
rect 5145 16294 5147 16346
rect 5327 16294 5329 16346
rect 5083 16292 5089 16294
rect 5145 16292 5169 16294
rect 5225 16292 5249 16294
rect 5305 16292 5329 16294
rect 5385 16292 5391 16294
rect 5083 16283 5391 16292
rect 12029 16348 12337 16357
rect 12029 16346 12035 16348
rect 12091 16346 12115 16348
rect 12171 16346 12195 16348
rect 12251 16346 12275 16348
rect 12331 16346 12337 16348
rect 12091 16294 12093 16346
rect 12273 16294 12275 16346
rect 12029 16292 12035 16294
rect 12091 16292 12115 16294
rect 12171 16292 12195 16294
rect 12251 16292 12275 16294
rect 12331 16292 12337 16294
rect 12029 16283 12337 16292
rect 4423 15804 4731 15813
rect 4423 15802 4429 15804
rect 4485 15802 4509 15804
rect 4565 15802 4589 15804
rect 4645 15802 4669 15804
rect 4725 15802 4731 15804
rect 4485 15750 4487 15802
rect 4667 15750 4669 15802
rect 4423 15748 4429 15750
rect 4485 15748 4509 15750
rect 4565 15748 4589 15750
rect 4645 15748 4669 15750
rect 4725 15748 4731 15750
rect 4423 15739 4731 15748
rect 11369 15804 11677 15813
rect 11369 15802 11375 15804
rect 11431 15802 11455 15804
rect 11511 15802 11535 15804
rect 11591 15802 11615 15804
rect 11671 15802 11677 15804
rect 11431 15750 11433 15802
rect 11613 15750 11615 15802
rect 11369 15748 11375 15750
rect 11431 15748 11455 15750
rect 11511 15748 11535 15750
rect 11591 15748 11615 15750
rect 11671 15748 11677 15750
rect 11369 15739 11677 15748
rect 5083 15260 5391 15269
rect 5083 15258 5089 15260
rect 5145 15258 5169 15260
rect 5225 15258 5249 15260
rect 5305 15258 5329 15260
rect 5385 15258 5391 15260
rect 5145 15206 5147 15258
rect 5327 15206 5329 15258
rect 5083 15204 5089 15206
rect 5145 15204 5169 15206
rect 5225 15204 5249 15206
rect 5305 15204 5329 15206
rect 5385 15204 5391 15206
rect 5083 15195 5391 15204
rect 12029 15260 12337 15269
rect 12029 15258 12035 15260
rect 12091 15258 12115 15260
rect 12171 15258 12195 15260
rect 12251 15258 12275 15260
rect 12331 15258 12337 15260
rect 12091 15206 12093 15258
rect 12273 15206 12275 15258
rect 12029 15204 12035 15206
rect 12091 15204 12115 15206
rect 12171 15204 12195 15206
rect 12251 15204 12275 15206
rect 12331 15204 12337 15206
rect 12029 15195 12337 15204
rect 4423 14716 4731 14725
rect 4423 14714 4429 14716
rect 4485 14714 4509 14716
rect 4565 14714 4589 14716
rect 4645 14714 4669 14716
rect 4725 14714 4731 14716
rect 4485 14662 4487 14714
rect 4667 14662 4669 14714
rect 4423 14660 4429 14662
rect 4485 14660 4509 14662
rect 4565 14660 4589 14662
rect 4645 14660 4669 14662
rect 4725 14660 4731 14662
rect 4423 14651 4731 14660
rect 11369 14716 11677 14725
rect 11369 14714 11375 14716
rect 11431 14714 11455 14716
rect 11511 14714 11535 14716
rect 11591 14714 11615 14716
rect 11671 14714 11677 14716
rect 11431 14662 11433 14714
rect 11613 14662 11615 14714
rect 11369 14660 11375 14662
rect 11431 14660 11455 14662
rect 11511 14660 11535 14662
rect 11591 14660 11615 14662
rect 11671 14660 11677 14662
rect 11369 14651 11677 14660
rect 5083 14172 5391 14181
rect 5083 14170 5089 14172
rect 5145 14170 5169 14172
rect 5225 14170 5249 14172
rect 5305 14170 5329 14172
rect 5385 14170 5391 14172
rect 5145 14118 5147 14170
rect 5327 14118 5329 14170
rect 5083 14116 5089 14118
rect 5145 14116 5169 14118
rect 5225 14116 5249 14118
rect 5305 14116 5329 14118
rect 5385 14116 5391 14118
rect 5083 14107 5391 14116
rect 12029 14172 12337 14181
rect 12029 14170 12035 14172
rect 12091 14170 12115 14172
rect 12171 14170 12195 14172
rect 12251 14170 12275 14172
rect 12331 14170 12337 14172
rect 12091 14118 12093 14170
rect 12273 14118 12275 14170
rect 12029 14116 12035 14118
rect 12091 14116 12115 14118
rect 12171 14116 12195 14118
rect 12251 14116 12275 14118
rect 12331 14116 12337 14118
rect 12029 14107 12337 14116
rect 4423 13628 4731 13637
rect 4423 13626 4429 13628
rect 4485 13626 4509 13628
rect 4565 13626 4589 13628
rect 4645 13626 4669 13628
rect 4725 13626 4731 13628
rect 4485 13574 4487 13626
rect 4667 13574 4669 13626
rect 4423 13572 4429 13574
rect 4485 13572 4509 13574
rect 4565 13572 4589 13574
rect 4645 13572 4669 13574
rect 4725 13572 4731 13574
rect 4423 13563 4731 13572
rect 11369 13628 11677 13637
rect 11369 13626 11375 13628
rect 11431 13626 11455 13628
rect 11511 13626 11535 13628
rect 11591 13626 11615 13628
rect 11671 13626 11677 13628
rect 11431 13574 11433 13626
rect 11613 13574 11615 13626
rect 11369 13572 11375 13574
rect 11431 13572 11455 13574
rect 11511 13572 11535 13574
rect 11591 13572 11615 13574
rect 11671 13572 11677 13574
rect 11369 13563 11677 13572
rect 5083 13084 5391 13093
rect 5083 13082 5089 13084
rect 5145 13082 5169 13084
rect 5225 13082 5249 13084
rect 5305 13082 5329 13084
rect 5385 13082 5391 13084
rect 5145 13030 5147 13082
rect 5327 13030 5329 13082
rect 5083 13028 5089 13030
rect 5145 13028 5169 13030
rect 5225 13028 5249 13030
rect 5305 13028 5329 13030
rect 5385 13028 5391 13030
rect 5083 13019 5391 13028
rect 12029 13084 12337 13093
rect 12029 13082 12035 13084
rect 12091 13082 12115 13084
rect 12171 13082 12195 13084
rect 12251 13082 12275 13084
rect 12331 13082 12337 13084
rect 12091 13030 12093 13082
rect 12273 13030 12275 13082
rect 12029 13028 12035 13030
rect 12091 13028 12115 13030
rect 12171 13028 12195 13030
rect 12251 13028 12275 13030
rect 12331 13028 12337 13030
rect 12029 13019 12337 13028
rect 4423 12540 4731 12549
rect 4423 12538 4429 12540
rect 4485 12538 4509 12540
rect 4565 12538 4589 12540
rect 4645 12538 4669 12540
rect 4725 12538 4731 12540
rect 4485 12486 4487 12538
rect 4667 12486 4669 12538
rect 4423 12484 4429 12486
rect 4485 12484 4509 12486
rect 4565 12484 4589 12486
rect 4645 12484 4669 12486
rect 4725 12484 4731 12486
rect 4423 12475 4731 12484
rect 11369 12540 11677 12549
rect 11369 12538 11375 12540
rect 11431 12538 11455 12540
rect 11511 12538 11535 12540
rect 11591 12538 11615 12540
rect 11671 12538 11677 12540
rect 11431 12486 11433 12538
rect 11613 12486 11615 12538
rect 11369 12484 11375 12486
rect 11431 12484 11455 12486
rect 11511 12484 11535 12486
rect 11591 12484 11615 12486
rect 11671 12484 11677 12486
rect 11369 12475 11677 12484
rect 5083 11996 5391 12005
rect 5083 11994 5089 11996
rect 5145 11994 5169 11996
rect 5225 11994 5249 11996
rect 5305 11994 5329 11996
rect 5385 11994 5391 11996
rect 5145 11942 5147 11994
rect 5327 11942 5329 11994
rect 5083 11940 5089 11942
rect 5145 11940 5169 11942
rect 5225 11940 5249 11942
rect 5305 11940 5329 11942
rect 5385 11940 5391 11942
rect 5083 11931 5391 11940
rect 12029 11996 12337 12005
rect 12029 11994 12035 11996
rect 12091 11994 12115 11996
rect 12171 11994 12195 11996
rect 12251 11994 12275 11996
rect 12331 11994 12337 11996
rect 12091 11942 12093 11994
rect 12273 11942 12275 11994
rect 12029 11940 12035 11942
rect 12091 11940 12115 11942
rect 12171 11940 12195 11942
rect 12251 11940 12275 11942
rect 12331 11940 12337 11942
rect 12029 11931 12337 11940
rect 4423 11452 4731 11461
rect 4423 11450 4429 11452
rect 4485 11450 4509 11452
rect 4565 11450 4589 11452
rect 4645 11450 4669 11452
rect 4725 11450 4731 11452
rect 4485 11398 4487 11450
rect 4667 11398 4669 11450
rect 4423 11396 4429 11398
rect 4485 11396 4509 11398
rect 4565 11396 4589 11398
rect 4645 11396 4669 11398
rect 4725 11396 4731 11398
rect 4423 11387 4731 11396
rect 11369 11452 11677 11461
rect 11369 11450 11375 11452
rect 11431 11450 11455 11452
rect 11511 11450 11535 11452
rect 11591 11450 11615 11452
rect 11671 11450 11677 11452
rect 11431 11398 11433 11450
rect 11613 11398 11615 11450
rect 11369 11396 11375 11398
rect 11431 11396 11455 11398
rect 11511 11396 11535 11398
rect 11591 11396 11615 11398
rect 11671 11396 11677 11398
rect 11369 11387 11677 11396
rect 13464 11218 13492 18702
rect 15856 12986 15884 27270
rect 16672 13320 16724 13326
rect 16672 13262 16724 13268
rect 16028 13184 16080 13190
rect 16028 13126 16080 13132
rect 16040 12986 16068 13126
rect 15844 12980 15896 12986
rect 15844 12922 15896 12928
rect 16028 12980 16080 12986
rect 16028 12922 16080 12928
rect 15476 12640 15528 12646
rect 15476 12582 15528 12588
rect 16304 12640 16356 12646
rect 16304 12582 16356 12588
rect 15488 12238 15516 12582
rect 16316 12306 16344 12582
rect 16304 12300 16356 12306
rect 16304 12242 16356 12248
rect 15476 12232 15528 12238
rect 15476 12174 15528 12180
rect 16488 12164 16540 12170
rect 16488 12106 16540 12112
rect 14924 12096 14976 12102
rect 14924 12038 14976 12044
rect 15108 12096 15160 12102
rect 15108 12038 15160 12044
rect 14936 11898 14964 12038
rect 14924 11892 14976 11898
rect 14924 11834 14976 11840
rect 15120 11558 15148 12038
rect 16500 11762 16528 12106
rect 16488 11756 16540 11762
rect 16488 11698 16540 11704
rect 14188 11552 14240 11558
rect 14188 11494 14240 11500
rect 15108 11552 15160 11558
rect 15108 11494 15160 11500
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 13820 11212 13872 11218
rect 13820 11154 13872 11160
rect 13544 11144 13596 11150
rect 13544 11086 13596 11092
rect 5083 10908 5391 10917
rect 5083 10906 5089 10908
rect 5145 10906 5169 10908
rect 5225 10906 5249 10908
rect 5305 10906 5329 10908
rect 5385 10906 5391 10908
rect 5145 10854 5147 10906
rect 5327 10854 5329 10906
rect 5083 10852 5089 10854
rect 5145 10852 5169 10854
rect 5225 10852 5249 10854
rect 5305 10852 5329 10854
rect 5385 10852 5391 10854
rect 5083 10843 5391 10852
rect 12029 10908 12337 10917
rect 12029 10906 12035 10908
rect 12091 10906 12115 10908
rect 12171 10906 12195 10908
rect 12251 10906 12275 10908
rect 12331 10906 12337 10908
rect 12091 10854 12093 10906
rect 12273 10854 12275 10906
rect 12029 10852 12035 10854
rect 12091 10852 12115 10854
rect 12171 10852 12195 10854
rect 12251 10852 12275 10854
rect 12331 10852 12337 10854
rect 12029 10843 12337 10852
rect 4423 10364 4731 10373
rect 4423 10362 4429 10364
rect 4485 10362 4509 10364
rect 4565 10362 4589 10364
rect 4645 10362 4669 10364
rect 4725 10362 4731 10364
rect 4485 10310 4487 10362
rect 4667 10310 4669 10362
rect 4423 10308 4429 10310
rect 4485 10308 4509 10310
rect 4565 10308 4589 10310
rect 4645 10308 4669 10310
rect 4725 10308 4731 10310
rect 4423 10299 4731 10308
rect 11369 10364 11677 10373
rect 11369 10362 11375 10364
rect 11431 10362 11455 10364
rect 11511 10362 11535 10364
rect 11591 10362 11615 10364
rect 11671 10362 11677 10364
rect 11431 10310 11433 10362
rect 11613 10310 11615 10362
rect 11369 10308 11375 10310
rect 11431 10308 11455 10310
rect 11511 10308 11535 10310
rect 11591 10308 11615 10310
rect 11671 10308 11677 10310
rect 11369 10299 11677 10308
rect 5083 9820 5391 9829
rect 5083 9818 5089 9820
rect 5145 9818 5169 9820
rect 5225 9818 5249 9820
rect 5305 9818 5329 9820
rect 5385 9818 5391 9820
rect 5145 9766 5147 9818
rect 5327 9766 5329 9818
rect 5083 9764 5089 9766
rect 5145 9764 5169 9766
rect 5225 9764 5249 9766
rect 5305 9764 5329 9766
rect 5385 9764 5391 9766
rect 5083 9755 5391 9764
rect 12029 9820 12337 9829
rect 12029 9818 12035 9820
rect 12091 9818 12115 9820
rect 12171 9818 12195 9820
rect 12251 9818 12275 9820
rect 12331 9818 12337 9820
rect 12091 9766 12093 9818
rect 12273 9766 12275 9818
rect 12029 9764 12035 9766
rect 12091 9764 12115 9766
rect 12171 9764 12195 9766
rect 12251 9764 12275 9766
rect 12331 9764 12337 9766
rect 12029 9755 12337 9764
rect 13556 9586 13584 11086
rect 13832 10810 13860 11154
rect 14200 11150 14228 11494
rect 15016 11212 15068 11218
rect 15016 11154 15068 11160
rect 14188 11144 14240 11150
rect 14188 11086 14240 11092
rect 15028 10810 15056 11154
rect 13820 10804 13872 10810
rect 13820 10746 13872 10752
rect 15016 10804 15068 10810
rect 15016 10746 15068 10752
rect 15016 10464 15068 10470
rect 15016 10406 15068 10412
rect 14372 9988 14424 9994
rect 14372 9930 14424 9936
rect 14384 9722 14412 9930
rect 14372 9716 14424 9722
rect 14372 9658 14424 9664
rect 13544 9580 13596 9586
rect 13544 9522 13596 9528
rect 4423 9276 4731 9285
rect 4423 9274 4429 9276
rect 4485 9274 4509 9276
rect 4565 9274 4589 9276
rect 4645 9274 4669 9276
rect 4725 9274 4731 9276
rect 4485 9222 4487 9274
rect 4667 9222 4669 9274
rect 4423 9220 4429 9222
rect 4485 9220 4509 9222
rect 4565 9220 4589 9222
rect 4645 9220 4669 9222
rect 4725 9220 4731 9222
rect 4423 9211 4731 9220
rect 11369 9276 11677 9285
rect 11369 9274 11375 9276
rect 11431 9274 11455 9276
rect 11511 9274 11535 9276
rect 11591 9274 11615 9276
rect 11671 9274 11677 9276
rect 11431 9222 11433 9274
rect 11613 9222 11615 9274
rect 11369 9220 11375 9222
rect 11431 9220 11455 9222
rect 11511 9220 11535 9222
rect 11591 9220 11615 9222
rect 11671 9220 11677 9222
rect 11369 9211 11677 9220
rect 940 8968 992 8974
rect 938 8936 940 8945
rect 992 8936 994 8945
rect 938 8871 994 8880
rect 5083 8732 5391 8741
rect 5083 8730 5089 8732
rect 5145 8730 5169 8732
rect 5225 8730 5249 8732
rect 5305 8730 5329 8732
rect 5385 8730 5391 8732
rect 5145 8678 5147 8730
rect 5327 8678 5329 8730
rect 5083 8676 5089 8678
rect 5145 8676 5169 8678
rect 5225 8676 5249 8678
rect 5305 8676 5329 8678
rect 5385 8676 5391 8678
rect 5083 8667 5391 8676
rect 12029 8732 12337 8741
rect 12029 8730 12035 8732
rect 12091 8730 12115 8732
rect 12171 8730 12195 8732
rect 12251 8730 12275 8732
rect 12331 8730 12337 8732
rect 12091 8678 12093 8730
rect 12273 8678 12275 8730
rect 12029 8676 12035 8678
rect 12091 8676 12115 8678
rect 12171 8676 12195 8678
rect 12251 8676 12275 8678
rect 12331 8676 12337 8678
rect 12029 8667 12337 8676
rect 4423 8188 4731 8197
rect 4423 8186 4429 8188
rect 4485 8186 4509 8188
rect 4565 8186 4589 8188
rect 4645 8186 4669 8188
rect 4725 8186 4731 8188
rect 4485 8134 4487 8186
rect 4667 8134 4669 8186
rect 4423 8132 4429 8134
rect 4485 8132 4509 8134
rect 4565 8132 4589 8134
rect 4645 8132 4669 8134
rect 4725 8132 4731 8134
rect 4423 8123 4731 8132
rect 11369 8188 11677 8197
rect 11369 8186 11375 8188
rect 11431 8186 11455 8188
rect 11511 8186 11535 8188
rect 11591 8186 11615 8188
rect 11671 8186 11677 8188
rect 11431 8134 11433 8186
rect 11613 8134 11615 8186
rect 11369 8132 11375 8134
rect 11431 8132 11455 8134
rect 11511 8132 11535 8134
rect 11591 8132 11615 8134
rect 11671 8132 11677 8134
rect 11369 8123 11677 8132
rect 5083 7644 5391 7653
rect 5083 7642 5089 7644
rect 5145 7642 5169 7644
rect 5225 7642 5249 7644
rect 5305 7642 5329 7644
rect 5385 7642 5391 7644
rect 5145 7590 5147 7642
rect 5327 7590 5329 7642
rect 5083 7588 5089 7590
rect 5145 7588 5169 7590
rect 5225 7588 5249 7590
rect 5305 7588 5329 7590
rect 5385 7588 5391 7590
rect 5083 7579 5391 7588
rect 12029 7644 12337 7653
rect 12029 7642 12035 7644
rect 12091 7642 12115 7644
rect 12171 7642 12195 7644
rect 12251 7642 12275 7644
rect 12331 7642 12337 7644
rect 12091 7590 12093 7642
rect 12273 7590 12275 7642
rect 12029 7588 12035 7590
rect 12091 7588 12115 7590
rect 12171 7588 12195 7590
rect 12251 7588 12275 7590
rect 12331 7588 12337 7590
rect 12029 7579 12337 7588
rect 4423 7100 4731 7109
rect 4423 7098 4429 7100
rect 4485 7098 4509 7100
rect 4565 7098 4589 7100
rect 4645 7098 4669 7100
rect 4725 7098 4731 7100
rect 4485 7046 4487 7098
rect 4667 7046 4669 7098
rect 4423 7044 4429 7046
rect 4485 7044 4509 7046
rect 4565 7044 4589 7046
rect 4645 7044 4669 7046
rect 4725 7044 4731 7046
rect 4423 7035 4731 7044
rect 11369 7100 11677 7109
rect 11369 7098 11375 7100
rect 11431 7098 11455 7100
rect 11511 7098 11535 7100
rect 11591 7098 11615 7100
rect 11671 7098 11677 7100
rect 11431 7046 11433 7098
rect 11613 7046 11615 7098
rect 11369 7044 11375 7046
rect 11431 7044 11455 7046
rect 11511 7044 11535 7046
rect 11591 7044 11615 7046
rect 11671 7044 11677 7046
rect 11369 7035 11677 7044
rect 5083 6556 5391 6565
rect 5083 6554 5089 6556
rect 5145 6554 5169 6556
rect 5225 6554 5249 6556
rect 5305 6554 5329 6556
rect 5385 6554 5391 6556
rect 5145 6502 5147 6554
rect 5327 6502 5329 6554
rect 5083 6500 5089 6502
rect 5145 6500 5169 6502
rect 5225 6500 5249 6502
rect 5305 6500 5329 6502
rect 5385 6500 5391 6502
rect 5083 6491 5391 6500
rect 12029 6556 12337 6565
rect 12029 6554 12035 6556
rect 12091 6554 12115 6556
rect 12171 6554 12195 6556
rect 12251 6554 12275 6556
rect 12331 6554 12337 6556
rect 12091 6502 12093 6554
rect 12273 6502 12275 6554
rect 12029 6500 12035 6502
rect 12091 6500 12115 6502
rect 12171 6500 12195 6502
rect 12251 6500 12275 6502
rect 12331 6500 12337 6502
rect 12029 6491 12337 6500
rect 4423 6012 4731 6021
rect 4423 6010 4429 6012
rect 4485 6010 4509 6012
rect 4565 6010 4589 6012
rect 4645 6010 4669 6012
rect 4725 6010 4731 6012
rect 4485 5958 4487 6010
rect 4667 5958 4669 6010
rect 4423 5956 4429 5958
rect 4485 5956 4509 5958
rect 4565 5956 4589 5958
rect 4645 5956 4669 5958
rect 4725 5956 4731 5958
rect 4423 5947 4731 5956
rect 11369 6012 11677 6021
rect 11369 6010 11375 6012
rect 11431 6010 11455 6012
rect 11511 6010 11535 6012
rect 11591 6010 11615 6012
rect 11671 6010 11677 6012
rect 11431 5958 11433 6010
rect 11613 5958 11615 6010
rect 11369 5956 11375 5958
rect 11431 5956 11455 5958
rect 11511 5956 11535 5958
rect 11591 5956 11615 5958
rect 11671 5956 11677 5958
rect 11369 5947 11677 5956
rect 5083 5468 5391 5477
rect 5083 5466 5089 5468
rect 5145 5466 5169 5468
rect 5225 5466 5249 5468
rect 5305 5466 5329 5468
rect 5385 5466 5391 5468
rect 5145 5414 5147 5466
rect 5327 5414 5329 5466
rect 5083 5412 5089 5414
rect 5145 5412 5169 5414
rect 5225 5412 5249 5414
rect 5305 5412 5329 5414
rect 5385 5412 5391 5414
rect 5083 5403 5391 5412
rect 12029 5468 12337 5477
rect 12029 5466 12035 5468
rect 12091 5466 12115 5468
rect 12171 5466 12195 5468
rect 12251 5466 12275 5468
rect 12331 5466 12337 5468
rect 12091 5414 12093 5466
rect 12273 5414 12275 5466
rect 12029 5412 12035 5414
rect 12091 5412 12115 5414
rect 12171 5412 12195 5414
rect 12251 5412 12275 5414
rect 12331 5412 12337 5414
rect 12029 5403 12337 5412
rect 4423 4924 4731 4933
rect 4423 4922 4429 4924
rect 4485 4922 4509 4924
rect 4565 4922 4589 4924
rect 4645 4922 4669 4924
rect 4725 4922 4731 4924
rect 4485 4870 4487 4922
rect 4667 4870 4669 4922
rect 4423 4868 4429 4870
rect 4485 4868 4509 4870
rect 4565 4868 4589 4870
rect 4645 4868 4669 4870
rect 4725 4868 4731 4870
rect 4423 4859 4731 4868
rect 11369 4924 11677 4933
rect 11369 4922 11375 4924
rect 11431 4922 11455 4924
rect 11511 4922 11535 4924
rect 11591 4922 11615 4924
rect 11671 4922 11677 4924
rect 11431 4870 11433 4922
rect 11613 4870 11615 4922
rect 11369 4868 11375 4870
rect 11431 4868 11455 4870
rect 11511 4868 11535 4870
rect 11591 4868 11615 4870
rect 11671 4868 11677 4870
rect 11369 4859 11677 4868
rect 5083 4380 5391 4389
rect 5083 4378 5089 4380
rect 5145 4378 5169 4380
rect 5225 4378 5249 4380
rect 5305 4378 5329 4380
rect 5385 4378 5391 4380
rect 5145 4326 5147 4378
rect 5327 4326 5329 4378
rect 5083 4324 5089 4326
rect 5145 4324 5169 4326
rect 5225 4324 5249 4326
rect 5305 4324 5329 4326
rect 5385 4324 5391 4326
rect 5083 4315 5391 4324
rect 12029 4380 12337 4389
rect 12029 4378 12035 4380
rect 12091 4378 12115 4380
rect 12171 4378 12195 4380
rect 12251 4378 12275 4380
rect 12331 4378 12337 4380
rect 12091 4326 12093 4378
rect 12273 4326 12275 4378
rect 12029 4324 12035 4326
rect 12091 4324 12115 4326
rect 12171 4324 12195 4326
rect 12251 4324 12275 4326
rect 12331 4324 12337 4326
rect 12029 4315 12337 4324
rect 4423 3836 4731 3845
rect 4423 3834 4429 3836
rect 4485 3834 4509 3836
rect 4565 3834 4589 3836
rect 4645 3834 4669 3836
rect 4725 3834 4731 3836
rect 4485 3782 4487 3834
rect 4667 3782 4669 3834
rect 4423 3780 4429 3782
rect 4485 3780 4509 3782
rect 4565 3780 4589 3782
rect 4645 3780 4669 3782
rect 4725 3780 4731 3782
rect 4423 3771 4731 3780
rect 11369 3836 11677 3845
rect 11369 3834 11375 3836
rect 11431 3834 11455 3836
rect 11511 3834 11535 3836
rect 11591 3834 11615 3836
rect 11671 3834 11677 3836
rect 11431 3782 11433 3834
rect 11613 3782 11615 3834
rect 11369 3780 11375 3782
rect 11431 3780 11455 3782
rect 11511 3780 11535 3782
rect 11591 3780 11615 3782
rect 11671 3780 11677 3782
rect 11369 3771 11677 3780
rect 5083 3292 5391 3301
rect 5083 3290 5089 3292
rect 5145 3290 5169 3292
rect 5225 3290 5249 3292
rect 5305 3290 5329 3292
rect 5385 3290 5391 3292
rect 5145 3238 5147 3290
rect 5327 3238 5329 3290
rect 5083 3236 5089 3238
rect 5145 3236 5169 3238
rect 5225 3236 5249 3238
rect 5305 3236 5329 3238
rect 5385 3236 5391 3238
rect 5083 3227 5391 3236
rect 12029 3292 12337 3301
rect 12029 3290 12035 3292
rect 12091 3290 12115 3292
rect 12171 3290 12195 3292
rect 12251 3290 12275 3292
rect 12331 3290 12337 3292
rect 12091 3238 12093 3290
rect 12273 3238 12275 3290
rect 12029 3236 12035 3238
rect 12091 3236 12115 3238
rect 12171 3236 12195 3238
rect 12251 3236 12275 3238
rect 12331 3236 12337 3238
rect 12029 3227 12337 3236
rect 4423 2748 4731 2757
rect 4423 2746 4429 2748
rect 4485 2746 4509 2748
rect 4565 2746 4589 2748
rect 4645 2746 4669 2748
rect 4725 2746 4731 2748
rect 4485 2694 4487 2746
rect 4667 2694 4669 2746
rect 4423 2692 4429 2694
rect 4485 2692 4509 2694
rect 4565 2692 4589 2694
rect 4645 2692 4669 2694
rect 4725 2692 4731 2694
rect 4423 2683 4731 2692
rect 11369 2748 11677 2757
rect 11369 2746 11375 2748
rect 11431 2746 11455 2748
rect 11511 2746 11535 2748
rect 11591 2746 11615 2748
rect 11671 2746 11677 2748
rect 11431 2694 11433 2746
rect 11613 2694 11615 2746
rect 11369 2692 11375 2694
rect 11431 2692 11455 2694
rect 11511 2692 11535 2694
rect 11591 2692 11615 2694
rect 11671 2692 11677 2694
rect 11369 2683 11677 2692
rect 13556 2514 13584 9522
rect 14740 9512 14792 9518
rect 15028 9500 15056 10406
rect 15120 10266 15148 11494
rect 16500 11218 16528 11698
rect 16684 11626 16712 13262
rect 17316 12776 17368 12782
rect 17316 12718 17368 12724
rect 17408 12776 17460 12782
rect 17408 12718 17460 12724
rect 17328 12646 17356 12718
rect 17316 12640 17368 12646
rect 17316 12582 17368 12588
rect 17328 11694 17356 12582
rect 17420 12102 17448 12718
rect 17604 12238 17632 27406
rect 20996 27396 21048 27402
rect 20996 27338 21048 27344
rect 18975 27228 19283 27237
rect 18975 27226 18981 27228
rect 19037 27226 19061 27228
rect 19117 27226 19141 27228
rect 19197 27226 19221 27228
rect 19277 27226 19283 27228
rect 19037 27174 19039 27226
rect 19219 27174 19221 27226
rect 18975 27172 18981 27174
rect 19037 27172 19061 27174
rect 19117 27172 19141 27174
rect 19197 27172 19221 27174
rect 19277 27172 19283 27174
rect 18975 27163 19283 27172
rect 18315 26684 18623 26693
rect 18315 26682 18321 26684
rect 18377 26682 18401 26684
rect 18457 26682 18481 26684
rect 18537 26682 18561 26684
rect 18617 26682 18623 26684
rect 18377 26630 18379 26682
rect 18559 26630 18561 26682
rect 18315 26628 18321 26630
rect 18377 26628 18401 26630
rect 18457 26628 18481 26630
rect 18537 26628 18561 26630
rect 18617 26628 18623 26630
rect 18315 26619 18623 26628
rect 18975 26140 19283 26149
rect 18975 26138 18981 26140
rect 19037 26138 19061 26140
rect 19117 26138 19141 26140
rect 19197 26138 19221 26140
rect 19277 26138 19283 26140
rect 19037 26086 19039 26138
rect 19219 26086 19221 26138
rect 18975 26084 18981 26086
rect 19037 26084 19061 26086
rect 19117 26084 19141 26086
rect 19197 26084 19221 26086
rect 19277 26084 19283 26086
rect 18975 26075 19283 26084
rect 18315 25596 18623 25605
rect 18315 25594 18321 25596
rect 18377 25594 18401 25596
rect 18457 25594 18481 25596
rect 18537 25594 18561 25596
rect 18617 25594 18623 25596
rect 18377 25542 18379 25594
rect 18559 25542 18561 25594
rect 18315 25540 18321 25542
rect 18377 25540 18401 25542
rect 18457 25540 18481 25542
rect 18537 25540 18561 25542
rect 18617 25540 18623 25542
rect 18315 25531 18623 25540
rect 18975 25052 19283 25061
rect 18975 25050 18981 25052
rect 19037 25050 19061 25052
rect 19117 25050 19141 25052
rect 19197 25050 19221 25052
rect 19277 25050 19283 25052
rect 19037 24998 19039 25050
rect 19219 24998 19221 25050
rect 18975 24996 18981 24998
rect 19037 24996 19061 24998
rect 19117 24996 19141 24998
rect 19197 24996 19221 24998
rect 19277 24996 19283 24998
rect 18975 24987 19283 24996
rect 18315 24508 18623 24517
rect 18315 24506 18321 24508
rect 18377 24506 18401 24508
rect 18457 24506 18481 24508
rect 18537 24506 18561 24508
rect 18617 24506 18623 24508
rect 18377 24454 18379 24506
rect 18559 24454 18561 24506
rect 18315 24452 18321 24454
rect 18377 24452 18401 24454
rect 18457 24452 18481 24454
rect 18537 24452 18561 24454
rect 18617 24452 18623 24454
rect 18315 24443 18623 24452
rect 18975 23964 19283 23973
rect 18975 23962 18981 23964
rect 19037 23962 19061 23964
rect 19117 23962 19141 23964
rect 19197 23962 19221 23964
rect 19277 23962 19283 23964
rect 19037 23910 19039 23962
rect 19219 23910 19221 23962
rect 18975 23908 18981 23910
rect 19037 23908 19061 23910
rect 19117 23908 19141 23910
rect 19197 23908 19221 23910
rect 19277 23908 19283 23910
rect 18975 23899 19283 23908
rect 18315 23420 18623 23429
rect 18315 23418 18321 23420
rect 18377 23418 18401 23420
rect 18457 23418 18481 23420
rect 18537 23418 18561 23420
rect 18617 23418 18623 23420
rect 18377 23366 18379 23418
rect 18559 23366 18561 23418
rect 18315 23364 18321 23366
rect 18377 23364 18401 23366
rect 18457 23364 18481 23366
rect 18537 23364 18561 23366
rect 18617 23364 18623 23366
rect 18315 23355 18623 23364
rect 18975 22876 19283 22885
rect 18975 22874 18981 22876
rect 19037 22874 19061 22876
rect 19117 22874 19141 22876
rect 19197 22874 19221 22876
rect 19277 22874 19283 22876
rect 19037 22822 19039 22874
rect 19219 22822 19221 22874
rect 18975 22820 18981 22822
rect 19037 22820 19061 22822
rect 19117 22820 19141 22822
rect 19197 22820 19221 22822
rect 19277 22820 19283 22822
rect 18975 22811 19283 22820
rect 18315 22332 18623 22341
rect 18315 22330 18321 22332
rect 18377 22330 18401 22332
rect 18457 22330 18481 22332
rect 18537 22330 18561 22332
rect 18617 22330 18623 22332
rect 18377 22278 18379 22330
rect 18559 22278 18561 22330
rect 18315 22276 18321 22278
rect 18377 22276 18401 22278
rect 18457 22276 18481 22278
rect 18537 22276 18561 22278
rect 18617 22276 18623 22278
rect 18315 22267 18623 22276
rect 18975 21788 19283 21797
rect 18975 21786 18981 21788
rect 19037 21786 19061 21788
rect 19117 21786 19141 21788
rect 19197 21786 19221 21788
rect 19277 21786 19283 21788
rect 19037 21734 19039 21786
rect 19219 21734 19221 21786
rect 18975 21732 18981 21734
rect 19037 21732 19061 21734
rect 19117 21732 19141 21734
rect 19197 21732 19221 21734
rect 19277 21732 19283 21734
rect 18975 21723 19283 21732
rect 18315 21244 18623 21253
rect 18315 21242 18321 21244
rect 18377 21242 18401 21244
rect 18457 21242 18481 21244
rect 18537 21242 18561 21244
rect 18617 21242 18623 21244
rect 18377 21190 18379 21242
rect 18559 21190 18561 21242
rect 18315 21188 18321 21190
rect 18377 21188 18401 21190
rect 18457 21188 18481 21190
rect 18537 21188 18561 21190
rect 18617 21188 18623 21190
rect 18315 21179 18623 21188
rect 18975 20700 19283 20709
rect 18975 20698 18981 20700
rect 19037 20698 19061 20700
rect 19117 20698 19141 20700
rect 19197 20698 19221 20700
rect 19277 20698 19283 20700
rect 19037 20646 19039 20698
rect 19219 20646 19221 20698
rect 18975 20644 18981 20646
rect 19037 20644 19061 20646
rect 19117 20644 19141 20646
rect 19197 20644 19221 20646
rect 19277 20644 19283 20646
rect 18975 20635 19283 20644
rect 18315 20156 18623 20165
rect 18315 20154 18321 20156
rect 18377 20154 18401 20156
rect 18457 20154 18481 20156
rect 18537 20154 18561 20156
rect 18617 20154 18623 20156
rect 18377 20102 18379 20154
rect 18559 20102 18561 20154
rect 18315 20100 18321 20102
rect 18377 20100 18401 20102
rect 18457 20100 18481 20102
rect 18537 20100 18561 20102
rect 18617 20100 18623 20102
rect 18315 20091 18623 20100
rect 18975 19612 19283 19621
rect 18975 19610 18981 19612
rect 19037 19610 19061 19612
rect 19117 19610 19141 19612
rect 19197 19610 19221 19612
rect 19277 19610 19283 19612
rect 19037 19558 19039 19610
rect 19219 19558 19221 19610
rect 18975 19556 18981 19558
rect 19037 19556 19061 19558
rect 19117 19556 19141 19558
rect 19197 19556 19221 19558
rect 19277 19556 19283 19558
rect 18975 19547 19283 19556
rect 18315 19068 18623 19077
rect 18315 19066 18321 19068
rect 18377 19066 18401 19068
rect 18457 19066 18481 19068
rect 18537 19066 18561 19068
rect 18617 19066 18623 19068
rect 18377 19014 18379 19066
rect 18559 19014 18561 19066
rect 18315 19012 18321 19014
rect 18377 19012 18401 19014
rect 18457 19012 18481 19014
rect 18537 19012 18561 19014
rect 18617 19012 18623 19014
rect 18315 19003 18623 19012
rect 18975 18524 19283 18533
rect 18975 18522 18981 18524
rect 19037 18522 19061 18524
rect 19117 18522 19141 18524
rect 19197 18522 19221 18524
rect 19277 18522 19283 18524
rect 19037 18470 19039 18522
rect 19219 18470 19221 18522
rect 18975 18468 18981 18470
rect 19037 18468 19061 18470
rect 19117 18468 19141 18470
rect 19197 18468 19221 18470
rect 19277 18468 19283 18470
rect 18975 18459 19283 18468
rect 18315 17980 18623 17989
rect 18315 17978 18321 17980
rect 18377 17978 18401 17980
rect 18457 17978 18481 17980
rect 18537 17978 18561 17980
rect 18617 17978 18623 17980
rect 18377 17926 18379 17978
rect 18559 17926 18561 17978
rect 18315 17924 18321 17926
rect 18377 17924 18401 17926
rect 18457 17924 18481 17926
rect 18537 17924 18561 17926
rect 18617 17924 18623 17926
rect 18315 17915 18623 17924
rect 18975 17436 19283 17445
rect 18975 17434 18981 17436
rect 19037 17434 19061 17436
rect 19117 17434 19141 17436
rect 19197 17434 19221 17436
rect 19277 17434 19283 17436
rect 19037 17382 19039 17434
rect 19219 17382 19221 17434
rect 18975 17380 18981 17382
rect 19037 17380 19061 17382
rect 19117 17380 19141 17382
rect 19197 17380 19221 17382
rect 19277 17380 19283 17382
rect 18975 17371 19283 17380
rect 18315 16892 18623 16901
rect 18315 16890 18321 16892
rect 18377 16890 18401 16892
rect 18457 16890 18481 16892
rect 18537 16890 18561 16892
rect 18617 16890 18623 16892
rect 18377 16838 18379 16890
rect 18559 16838 18561 16890
rect 18315 16836 18321 16838
rect 18377 16836 18401 16838
rect 18457 16836 18481 16838
rect 18537 16836 18561 16838
rect 18617 16836 18623 16838
rect 18315 16827 18623 16836
rect 18975 16348 19283 16357
rect 18975 16346 18981 16348
rect 19037 16346 19061 16348
rect 19117 16346 19141 16348
rect 19197 16346 19221 16348
rect 19277 16346 19283 16348
rect 19037 16294 19039 16346
rect 19219 16294 19221 16346
rect 18975 16292 18981 16294
rect 19037 16292 19061 16294
rect 19117 16292 19141 16294
rect 19197 16292 19221 16294
rect 19277 16292 19283 16294
rect 18975 16283 19283 16292
rect 18315 15804 18623 15813
rect 18315 15802 18321 15804
rect 18377 15802 18401 15804
rect 18457 15802 18481 15804
rect 18537 15802 18561 15804
rect 18617 15802 18623 15804
rect 18377 15750 18379 15802
rect 18559 15750 18561 15802
rect 18315 15748 18321 15750
rect 18377 15748 18401 15750
rect 18457 15748 18481 15750
rect 18537 15748 18561 15750
rect 18617 15748 18623 15750
rect 18315 15739 18623 15748
rect 18975 15260 19283 15269
rect 18975 15258 18981 15260
rect 19037 15258 19061 15260
rect 19117 15258 19141 15260
rect 19197 15258 19221 15260
rect 19277 15258 19283 15260
rect 19037 15206 19039 15258
rect 19219 15206 19221 15258
rect 18975 15204 18981 15206
rect 19037 15204 19061 15206
rect 19117 15204 19141 15206
rect 19197 15204 19221 15206
rect 19277 15204 19283 15206
rect 18975 15195 19283 15204
rect 18315 14716 18623 14725
rect 18315 14714 18321 14716
rect 18377 14714 18401 14716
rect 18457 14714 18481 14716
rect 18537 14714 18561 14716
rect 18617 14714 18623 14716
rect 18377 14662 18379 14714
rect 18559 14662 18561 14714
rect 18315 14660 18321 14662
rect 18377 14660 18401 14662
rect 18457 14660 18481 14662
rect 18537 14660 18561 14662
rect 18617 14660 18623 14662
rect 18315 14651 18623 14660
rect 18975 14172 19283 14181
rect 18975 14170 18981 14172
rect 19037 14170 19061 14172
rect 19117 14170 19141 14172
rect 19197 14170 19221 14172
rect 19277 14170 19283 14172
rect 19037 14118 19039 14170
rect 19219 14118 19221 14170
rect 18975 14116 18981 14118
rect 19037 14116 19061 14118
rect 19117 14116 19141 14118
rect 19197 14116 19221 14118
rect 19277 14116 19283 14118
rect 18975 14107 19283 14116
rect 18315 13628 18623 13637
rect 18315 13626 18321 13628
rect 18377 13626 18401 13628
rect 18457 13626 18481 13628
rect 18537 13626 18561 13628
rect 18617 13626 18623 13628
rect 18377 13574 18379 13626
rect 18559 13574 18561 13626
rect 18315 13572 18321 13574
rect 18377 13572 18401 13574
rect 18457 13572 18481 13574
rect 18537 13572 18561 13574
rect 18617 13572 18623 13574
rect 18315 13563 18623 13572
rect 18975 13084 19283 13093
rect 18975 13082 18981 13084
rect 19037 13082 19061 13084
rect 19117 13082 19141 13084
rect 19197 13082 19221 13084
rect 19277 13082 19283 13084
rect 19037 13030 19039 13082
rect 19219 13030 19221 13082
rect 18975 13028 18981 13030
rect 19037 13028 19061 13030
rect 19117 13028 19141 13030
rect 19197 13028 19221 13030
rect 19277 13028 19283 13030
rect 18975 13019 19283 13028
rect 19248 12844 19300 12850
rect 19248 12786 19300 12792
rect 18880 12708 18932 12714
rect 18880 12650 18932 12656
rect 18315 12540 18623 12549
rect 18315 12538 18321 12540
rect 18377 12538 18401 12540
rect 18457 12538 18481 12540
rect 18537 12538 18561 12540
rect 18617 12538 18623 12540
rect 18377 12486 18379 12538
rect 18559 12486 18561 12538
rect 18315 12484 18321 12486
rect 18377 12484 18401 12486
rect 18457 12484 18481 12486
rect 18537 12484 18561 12486
rect 18617 12484 18623 12486
rect 18315 12475 18623 12484
rect 17960 12300 18012 12306
rect 17960 12242 18012 12248
rect 17592 12232 17644 12238
rect 17592 12174 17644 12180
rect 17408 12096 17460 12102
rect 17408 12038 17460 12044
rect 17316 11688 17368 11694
rect 17316 11630 17368 11636
rect 16672 11620 16724 11626
rect 16672 11562 16724 11568
rect 17224 11552 17276 11558
rect 17224 11494 17276 11500
rect 16580 11348 16632 11354
rect 16580 11290 16632 11296
rect 16488 11212 16540 11218
rect 16488 11154 16540 11160
rect 15752 11076 15804 11082
rect 15752 11018 15804 11024
rect 15108 10260 15160 10266
rect 15108 10202 15160 10208
rect 14792 9472 15056 9500
rect 14740 9454 14792 9460
rect 14740 9376 14792 9382
rect 14740 9318 14792 9324
rect 14752 8906 14780 9318
rect 15028 9042 15056 9472
rect 15016 9036 15068 9042
rect 15016 8978 15068 8984
rect 14740 8900 14792 8906
rect 14740 8842 14792 8848
rect 14096 8832 14148 8838
rect 14096 8774 14148 8780
rect 14108 8566 14136 8774
rect 15120 8634 15148 10202
rect 15764 10062 15792 11018
rect 15936 11008 15988 11014
rect 15936 10950 15988 10956
rect 16304 11008 16356 11014
rect 16304 10950 16356 10956
rect 15948 10606 15976 10950
rect 15936 10600 15988 10606
rect 15936 10542 15988 10548
rect 16316 10266 16344 10950
rect 16396 10668 16448 10674
rect 16396 10610 16448 10616
rect 16304 10260 16356 10266
rect 16304 10202 16356 10208
rect 15752 10056 15804 10062
rect 15752 9998 15804 10004
rect 15108 8628 15160 8634
rect 15108 8570 15160 8576
rect 14096 8560 14148 8566
rect 14096 8502 14148 8508
rect 15120 8090 15148 8570
rect 15764 8566 15792 9998
rect 15936 9920 15988 9926
rect 15936 9862 15988 9868
rect 15948 9722 15976 9862
rect 15936 9716 15988 9722
rect 15936 9658 15988 9664
rect 16408 9518 16436 10610
rect 16592 10606 16620 11290
rect 17236 10810 17264 11494
rect 17316 11008 17368 11014
rect 17316 10950 17368 10956
rect 17328 10810 17356 10950
rect 17224 10804 17276 10810
rect 17224 10746 17276 10752
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 16488 10600 16540 10606
rect 16488 10542 16540 10548
rect 16580 10600 16632 10606
rect 16580 10542 16632 10548
rect 16500 9518 16528 10542
rect 17420 9674 17448 12038
rect 17604 11898 17632 12174
rect 17592 11892 17644 11898
rect 17592 11834 17644 11840
rect 17776 11688 17828 11694
rect 17776 11630 17828 11636
rect 17500 11552 17552 11558
rect 17500 11494 17552 11500
rect 17052 9646 17448 9674
rect 16396 9512 16448 9518
rect 16396 9454 16448 9460
rect 16488 9512 16540 9518
rect 16488 9454 16540 9460
rect 16764 9376 16816 9382
rect 16764 9318 16816 9324
rect 16776 9081 16804 9318
rect 17052 9110 17080 9646
rect 17408 9580 17460 9586
rect 17328 9540 17408 9568
rect 17328 9382 17356 9540
rect 17408 9522 17460 9528
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 17316 9376 17368 9382
rect 17316 9318 17368 9324
rect 17040 9104 17092 9110
rect 16762 9072 16818 9081
rect 15936 9036 15988 9042
rect 17040 9046 17092 9052
rect 16762 9007 16818 9016
rect 17132 9036 17184 9042
rect 15936 8978 15988 8984
rect 17132 8978 17184 8984
rect 15948 8634 15976 8978
rect 16028 8968 16080 8974
rect 16028 8910 16080 8916
rect 16396 8968 16448 8974
rect 16396 8910 16448 8916
rect 16040 8634 16068 8910
rect 16212 8832 16264 8838
rect 16212 8774 16264 8780
rect 15936 8628 15988 8634
rect 15936 8570 15988 8576
rect 16028 8628 16080 8634
rect 16028 8570 16080 8576
rect 15752 8560 15804 8566
rect 15752 8502 15804 8508
rect 15108 8084 15160 8090
rect 15108 8026 15160 8032
rect 15764 7478 15792 8502
rect 16224 7478 16252 8774
rect 16408 8430 16436 8910
rect 16396 8424 16448 8430
rect 16396 8366 16448 8372
rect 16408 7546 16436 8366
rect 17144 8090 17172 8978
rect 17236 8566 17264 9318
rect 17512 9042 17540 11494
rect 17788 11218 17816 11630
rect 17776 11212 17828 11218
rect 17776 11154 17828 11160
rect 17788 10606 17816 11154
rect 17972 10674 18000 12242
rect 18892 11778 18920 12650
rect 19260 12374 19288 12786
rect 19248 12368 19300 12374
rect 19248 12310 19300 12316
rect 18975 11996 19283 12005
rect 18975 11994 18981 11996
rect 19037 11994 19061 11996
rect 19117 11994 19141 11996
rect 19197 11994 19221 11996
rect 19277 11994 19283 11996
rect 19037 11942 19039 11994
rect 19219 11942 19221 11994
rect 18975 11940 18981 11942
rect 19037 11940 19061 11942
rect 19117 11940 19141 11942
rect 19197 11940 19221 11942
rect 19277 11940 19283 11942
rect 18975 11931 19283 11940
rect 18892 11762 19012 11778
rect 18892 11756 19024 11762
rect 18892 11750 18972 11756
rect 18972 11698 19024 11704
rect 19248 11756 19300 11762
rect 19248 11698 19300 11704
rect 18236 11620 18288 11626
rect 18236 11562 18288 11568
rect 18052 11552 18104 11558
rect 18052 11494 18104 11500
rect 18064 11286 18092 11494
rect 18052 11280 18104 11286
rect 18052 11222 18104 11228
rect 17960 10668 18012 10674
rect 17960 10610 18012 10616
rect 17776 10600 17828 10606
rect 17776 10542 17828 10548
rect 17592 9920 17644 9926
rect 17592 9862 17644 9868
rect 17604 9674 17632 9862
rect 17604 9646 17705 9674
rect 17677 9518 17705 9646
rect 17677 9512 17736 9518
rect 17677 9472 17684 9512
rect 17788 9489 17816 10542
rect 17972 9674 18000 10610
rect 18064 9674 18092 11222
rect 18144 11008 18196 11014
rect 18144 10950 18196 10956
rect 18156 10810 18184 10950
rect 18144 10804 18196 10810
rect 18144 10746 18196 10752
rect 18248 10606 18276 11562
rect 18315 11452 18623 11461
rect 18315 11450 18321 11452
rect 18377 11450 18401 11452
rect 18457 11450 18481 11452
rect 18537 11450 18561 11452
rect 18617 11450 18623 11452
rect 18377 11398 18379 11450
rect 18559 11398 18561 11450
rect 18315 11396 18321 11398
rect 18377 11396 18401 11398
rect 18457 11396 18481 11398
rect 18537 11396 18561 11398
rect 18617 11396 18623 11398
rect 18315 11387 18623 11396
rect 19260 11354 19288 11698
rect 19984 11688 20036 11694
rect 19984 11630 20036 11636
rect 20168 11688 20220 11694
rect 20168 11630 20220 11636
rect 19340 11620 19392 11626
rect 19340 11562 19392 11568
rect 19248 11348 19300 11354
rect 19248 11290 19300 11296
rect 19352 11150 19380 11562
rect 19432 11552 19484 11558
rect 19432 11494 19484 11500
rect 18788 11144 18840 11150
rect 18788 11086 18840 11092
rect 19340 11144 19392 11150
rect 19340 11086 19392 11092
rect 18236 10600 18288 10606
rect 18236 10542 18288 10548
rect 18236 10464 18288 10470
rect 18236 10406 18288 10412
rect 18696 10464 18748 10470
rect 18696 10406 18748 10412
rect 18248 10198 18276 10406
rect 18315 10364 18623 10373
rect 18315 10362 18321 10364
rect 18377 10362 18401 10364
rect 18457 10362 18481 10364
rect 18537 10362 18561 10364
rect 18617 10362 18623 10364
rect 18377 10310 18379 10362
rect 18559 10310 18561 10362
rect 18315 10308 18321 10310
rect 18377 10308 18401 10310
rect 18457 10308 18481 10310
rect 18537 10308 18561 10310
rect 18617 10308 18623 10310
rect 18315 10299 18623 10308
rect 18708 10266 18736 10406
rect 18800 10266 18828 11086
rect 18880 11008 18932 11014
rect 18880 10950 18932 10956
rect 18696 10260 18748 10266
rect 18696 10202 18748 10208
rect 18788 10260 18840 10266
rect 18788 10202 18840 10208
rect 18236 10192 18288 10198
rect 18236 10134 18288 10140
rect 18696 9988 18748 9994
rect 18696 9930 18748 9936
rect 17972 9646 18026 9674
rect 18064 9646 18276 9674
rect 17684 9454 17736 9460
rect 17774 9480 17830 9489
rect 17774 9415 17830 9424
rect 17998 9432 18026 9646
rect 18248 9586 18276 9646
rect 18236 9580 18288 9586
rect 18236 9522 18288 9528
rect 18144 9444 18196 9450
rect 17998 9404 18092 9432
rect 17684 9376 17736 9382
rect 17684 9318 17736 9324
rect 17774 9344 17830 9353
rect 17696 9042 17724 9318
rect 17774 9279 17830 9288
rect 17788 9178 17816 9279
rect 17776 9172 17828 9178
rect 17776 9114 17828 9120
rect 17500 9036 17552 9042
rect 17500 8978 17552 8984
rect 17684 9036 17736 9042
rect 17684 8978 17736 8984
rect 17224 8560 17276 8566
rect 17224 8502 17276 8508
rect 17132 8084 17184 8090
rect 17132 8026 17184 8032
rect 17040 7744 17092 7750
rect 17040 7686 17092 7692
rect 16396 7540 16448 7546
rect 16396 7482 16448 7488
rect 15752 7472 15804 7478
rect 15752 7414 15804 7420
rect 16212 7472 16264 7478
rect 16212 7414 16264 7420
rect 16580 7336 16632 7342
rect 16580 7278 16632 7284
rect 16592 6662 16620 7278
rect 17052 7002 17080 7686
rect 17040 6996 17092 7002
rect 17040 6938 17092 6944
rect 16580 6656 16632 6662
rect 16580 6598 16632 6604
rect 16592 6254 16620 6598
rect 16580 6248 16632 6254
rect 16580 6190 16632 6196
rect 16592 5574 16620 6190
rect 16580 5568 16632 5574
rect 16580 5510 16632 5516
rect 16592 5166 16620 5510
rect 16580 5160 16632 5166
rect 16580 5102 16632 5108
rect 16592 4690 16620 5102
rect 16580 4684 16632 4690
rect 16580 4626 16632 4632
rect 16120 4548 16172 4554
rect 16120 4490 16172 4496
rect 16132 4282 16160 4490
rect 16120 4276 16172 4282
rect 16120 4218 16172 4224
rect 16592 3602 16620 4626
rect 17130 4176 17186 4185
rect 17130 4111 17132 4120
rect 17184 4111 17186 4120
rect 17132 4082 17184 4088
rect 16580 3596 16632 3602
rect 16580 3538 16632 3544
rect 16856 3460 16908 3466
rect 16856 3402 16908 3408
rect 16868 3194 16896 3402
rect 16856 3188 16908 3194
rect 16856 3130 16908 3136
rect 17236 2774 17264 8502
rect 17500 8084 17552 8090
rect 17500 8026 17552 8032
rect 17512 7546 17540 8026
rect 17696 7970 17724 8978
rect 17788 8498 17816 9114
rect 17776 8492 17828 8498
rect 17776 8434 17828 8440
rect 17604 7942 17724 7970
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 17604 7410 17632 7942
rect 17684 7880 17736 7886
rect 17776 7880 17828 7886
rect 17684 7822 17736 7828
rect 17774 7848 17776 7857
rect 17828 7848 17830 7857
rect 17696 7546 17724 7822
rect 17774 7783 17830 7792
rect 17684 7540 17736 7546
rect 17684 7482 17736 7488
rect 17592 7404 17644 7410
rect 17592 7346 17644 7352
rect 17604 6984 17632 7346
rect 17880 7313 17908 7958
rect 17866 7304 17922 7313
rect 17866 7239 17922 7248
rect 17684 6996 17736 7002
rect 17604 6956 17684 6984
rect 17684 6938 17736 6944
rect 17408 6248 17460 6254
rect 17408 6190 17460 6196
rect 17420 4826 17448 6190
rect 17880 5710 17908 7239
rect 18064 5930 18092 9404
rect 18144 9386 18196 9392
rect 18156 8566 18184 9386
rect 18236 9376 18288 9382
rect 18236 9318 18288 9324
rect 18248 8956 18276 9318
rect 18315 9276 18623 9285
rect 18315 9274 18321 9276
rect 18377 9274 18401 9276
rect 18457 9274 18481 9276
rect 18537 9274 18561 9276
rect 18617 9274 18623 9276
rect 18377 9222 18379 9274
rect 18559 9222 18561 9274
rect 18315 9220 18321 9222
rect 18377 9220 18401 9222
rect 18457 9220 18481 9222
rect 18537 9220 18561 9222
rect 18617 9220 18623 9222
rect 18315 9211 18623 9220
rect 18604 8968 18656 8974
rect 18248 8928 18604 8956
rect 18604 8910 18656 8916
rect 18236 8832 18288 8838
rect 18236 8774 18288 8780
rect 18144 8560 18196 8566
rect 18144 8502 18196 8508
rect 18248 7886 18276 8774
rect 18616 8378 18644 8910
rect 18708 8566 18736 9930
rect 18800 9586 18828 10202
rect 18892 9994 18920 10950
rect 18975 10908 19283 10917
rect 18975 10906 18981 10908
rect 19037 10906 19061 10908
rect 19117 10906 19141 10908
rect 19197 10906 19221 10908
rect 19277 10906 19283 10908
rect 19037 10854 19039 10906
rect 19219 10854 19221 10906
rect 18975 10852 18981 10854
rect 19037 10852 19061 10854
rect 19117 10852 19141 10854
rect 19197 10852 19221 10854
rect 19277 10852 19283 10854
rect 18975 10843 19283 10852
rect 19444 10606 19472 11494
rect 19708 10736 19760 10742
rect 19708 10678 19760 10684
rect 19432 10600 19484 10606
rect 19432 10542 19484 10548
rect 18880 9988 18932 9994
rect 18880 9930 18932 9936
rect 19616 9988 19668 9994
rect 19616 9930 19668 9936
rect 18975 9820 19283 9829
rect 18975 9818 18981 9820
rect 19037 9818 19061 9820
rect 19117 9818 19141 9820
rect 19197 9818 19221 9820
rect 19277 9818 19283 9820
rect 19037 9766 19039 9818
rect 19219 9766 19221 9818
rect 18975 9764 18981 9766
rect 19037 9764 19061 9766
rect 19117 9764 19141 9766
rect 19197 9764 19221 9766
rect 19277 9764 19283 9766
rect 18975 9755 19283 9764
rect 19628 9722 19656 9930
rect 19616 9716 19668 9722
rect 19616 9658 19668 9664
rect 18788 9580 18840 9586
rect 18788 9522 18840 9528
rect 18788 9444 18840 9450
rect 18788 9386 18840 9392
rect 19432 9444 19484 9450
rect 19432 9386 19484 9392
rect 18696 8560 18748 8566
rect 18696 8502 18748 8508
rect 18616 8350 18736 8378
rect 18315 8188 18623 8197
rect 18315 8186 18321 8188
rect 18377 8186 18401 8188
rect 18457 8186 18481 8188
rect 18537 8186 18561 8188
rect 18617 8186 18623 8188
rect 18377 8134 18379 8186
rect 18559 8134 18561 8186
rect 18315 8132 18321 8134
rect 18377 8132 18401 8134
rect 18457 8132 18481 8134
rect 18537 8132 18561 8134
rect 18617 8132 18623 8134
rect 18315 8123 18623 8132
rect 18708 8090 18736 8350
rect 18696 8084 18748 8090
rect 18696 8026 18748 8032
rect 18328 8016 18380 8022
rect 18328 7958 18380 7964
rect 18236 7880 18288 7886
rect 18236 7822 18288 7828
rect 18236 7744 18288 7750
rect 18236 7686 18288 7692
rect 18248 6798 18276 7686
rect 18340 7546 18368 7958
rect 18696 7880 18748 7886
rect 18694 7848 18696 7857
rect 18748 7848 18750 7857
rect 18694 7783 18750 7792
rect 18708 7546 18736 7783
rect 18328 7540 18380 7546
rect 18328 7482 18380 7488
rect 18696 7540 18748 7546
rect 18696 7482 18748 7488
rect 18696 7336 18748 7342
rect 18696 7278 18748 7284
rect 18315 7100 18623 7109
rect 18315 7098 18321 7100
rect 18377 7098 18401 7100
rect 18457 7098 18481 7100
rect 18537 7098 18561 7100
rect 18617 7098 18623 7100
rect 18377 7046 18379 7098
rect 18559 7046 18561 7098
rect 18315 7044 18321 7046
rect 18377 7044 18401 7046
rect 18457 7044 18481 7046
rect 18537 7044 18561 7046
rect 18617 7044 18623 7046
rect 18315 7035 18623 7044
rect 18708 7002 18736 7278
rect 18696 6996 18748 7002
rect 18696 6938 18748 6944
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 18696 6792 18748 6798
rect 18696 6734 18748 6740
rect 18800 6746 18828 9386
rect 19248 9376 19300 9382
rect 19248 9318 19300 9324
rect 19340 9376 19392 9382
rect 19340 9318 19392 9324
rect 19260 9178 19288 9318
rect 19248 9172 19300 9178
rect 19248 9114 19300 9120
rect 18878 9072 18934 9081
rect 18878 9007 18880 9016
rect 18932 9007 18934 9016
rect 18880 8978 18932 8984
rect 19352 8838 19380 9318
rect 19444 9110 19472 9386
rect 19432 9104 19484 9110
rect 19432 9046 19484 9052
rect 19340 8832 19392 8838
rect 19340 8774 19392 8780
rect 18975 8732 19283 8741
rect 18975 8730 18981 8732
rect 19037 8730 19061 8732
rect 19117 8730 19141 8732
rect 19197 8730 19221 8732
rect 19277 8730 19283 8732
rect 19037 8678 19039 8730
rect 19219 8678 19221 8730
rect 18975 8676 18981 8678
rect 19037 8676 19061 8678
rect 19117 8676 19141 8678
rect 19197 8676 19221 8678
rect 19277 8676 19283 8678
rect 18975 8667 19283 8676
rect 19352 8634 19380 8774
rect 19340 8628 19392 8634
rect 19340 8570 19392 8576
rect 19444 7886 19472 9046
rect 19432 7880 19484 7886
rect 19432 7822 19484 7828
rect 18975 7644 19283 7653
rect 18975 7642 18981 7644
rect 19037 7642 19061 7644
rect 19117 7642 19141 7644
rect 19197 7642 19221 7644
rect 19277 7642 19283 7644
rect 19037 7590 19039 7642
rect 19219 7590 19221 7642
rect 18975 7588 18981 7590
rect 19037 7588 19061 7590
rect 19117 7588 19141 7590
rect 19197 7588 19221 7590
rect 19277 7588 19283 7590
rect 18975 7579 19283 7588
rect 19720 7478 19748 10678
rect 19996 10470 20024 11630
rect 19984 10464 20036 10470
rect 19984 10406 20036 10412
rect 19996 8498 20024 10406
rect 20076 9512 20128 9518
rect 20076 9454 20128 9460
rect 19984 8492 20036 8498
rect 19984 8434 20036 8440
rect 20088 7886 20116 9454
rect 20180 9450 20208 11630
rect 21008 11354 21036 27338
rect 21652 11558 21680 27542
rect 25148 27538 25176 29200
rect 25261 27772 25569 27781
rect 25261 27770 25267 27772
rect 25323 27770 25347 27772
rect 25403 27770 25427 27772
rect 25483 27770 25507 27772
rect 25563 27770 25569 27772
rect 25323 27718 25325 27770
rect 25505 27718 25507 27770
rect 25261 27716 25267 27718
rect 25323 27716 25347 27718
rect 25403 27716 25427 27718
rect 25483 27716 25507 27718
rect 25563 27716 25569 27718
rect 25261 27707 25569 27716
rect 25136 27532 25188 27538
rect 25136 27474 25188 27480
rect 25921 27228 26229 27237
rect 25921 27226 25927 27228
rect 25983 27226 26007 27228
rect 26063 27226 26087 27228
rect 26143 27226 26167 27228
rect 26223 27226 26229 27228
rect 25983 27174 25985 27226
rect 26165 27174 26167 27226
rect 25921 27172 25927 27174
rect 25983 27172 26007 27174
rect 26063 27172 26087 27174
rect 26143 27172 26167 27174
rect 26223 27172 26229 27174
rect 25921 27163 26229 27172
rect 25261 26684 25569 26693
rect 25261 26682 25267 26684
rect 25323 26682 25347 26684
rect 25403 26682 25427 26684
rect 25483 26682 25507 26684
rect 25563 26682 25569 26684
rect 25323 26630 25325 26682
rect 25505 26630 25507 26682
rect 25261 26628 25267 26630
rect 25323 26628 25347 26630
rect 25403 26628 25427 26630
rect 25483 26628 25507 26630
rect 25563 26628 25569 26630
rect 25261 26619 25569 26628
rect 25921 26140 26229 26149
rect 25921 26138 25927 26140
rect 25983 26138 26007 26140
rect 26063 26138 26087 26140
rect 26143 26138 26167 26140
rect 26223 26138 26229 26140
rect 25983 26086 25985 26138
rect 26165 26086 26167 26138
rect 25921 26084 25927 26086
rect 25983 26084 26007 26086
rect 26063 26084 26087 26086
rect 26143 26084 26167 26086
rect 26223 26084 26229 26086
rect 25921 26075 26229 26084
rect 25261 25596 25569 25605
rect 25261 25594 25267 25596
rect 25323 25594 25347 25596
rect 25403 25594 25427 25596
rect 25483 25594 25507 25596
rect 25563 25594 25569 25596
rect 25323 25542 25325 25594
rect 25505 25542 25507 25594
rect 25261 25540 25267 25542
rect 25323 25540 25347 25542
rect 25403 25540 25427 25542
rect 25483 25540 25507 25542
rect 25563 25540 25569 25542
rect 25261 25531 25569 25540
rect 28264 25288 28316 25294
rect 28540 25288 28592 25294
rect 28264 25230 28316 25236
rect 28538 25256 28540 25265
rect 28592 25256 28594 25265
rect 25921 25052 26229 25061
rect 25921 25050 25927 25052
rect 25983 25050 26007 25052
rect 26063 25050 26087 25052
rect 26143 25050 26167 25052
rect 26223 25050 26229 25052
rect 25983 24998 25985 25050
rect 26165 24998 26167 25050
rect 25921 24996 25927 24998
rect 25983 24996 26007 24998
rect 26063 24996 26087 24998
rect 26143 24996 26167 24998
rect 26223 24996 26229 24998
rect 25921 24987 26229 24996
rect 25261 24508 25569 24517
rect 25261 24506 25267 24508
rect 25323 24506 25347 24508
rect 25403 24506 25427 24508
rect 25483 24506 25507 24508
rect 25563 24506 25569 24508
rect 25323 24454 25325 24506
rect 25505 24454 25507 24506
rect 25261 24452 25267 24454
rect 25323 24452 25347 24454
rect 25403 24452 25427 24454
rect 25483 24452 25507 24454
rect 25563 24452 25569 24454
rect 25261 24443 25569 24452
rect 25921 23964 26229 23973
rect 25921 23962 25927 23964
rect 25983 23962 26007 23964
rect 26063 23962 26087 23964
rect 26143 23962 26167 23964
rect 26223 23962 26229 23964
rect 25983 23910 25985 23962
rect 26165 23910 26167 23962
rect 25921 23908 25927 23910
rect 25983 23908 26007 23910
rect 26063 23908 26087 23910
rect 26143 23908 26167 23910
rect 26223 23908 26229 23910
rect 25921 23899 26229 23908
rect 25261 23420 25569 23429
rect 25261 23418 25267 23420
rect 25323 23418 25347 23420
rect 25403 23418 25427 23420
rect 25483 23418 25507 23420
rect 25563 23418 25569 23420
rect 25323 23366 25325 23418
rect 25505 23366 25507 23418
rect 25261 23364 25267 23366
rect 25323 23364 25347 23366
rect 25403 23364 25427 23366
rect 25483 23364 25507 23366
rect 25563 23364 25569 23366
rect 25261 23355 25569 23364
rect 25921 22876 26229 22885
rect 25921 22874 25927 22876
rect 25983 22874 26007 22876
rect 26063 22874 26087 22876
rect 26143 22874 26167 22876
rect 26223 22874 26229 22876
rect 25983 22822 25985 22874
rect 26165 22822 26167 22874
rect 25921 22820 25927 22822
rect 25983 22820 26007 22822
rect 26063 22820 26087 22822
rect 26143 22820 26167 22822
rect 26223 22820 26229 22822
rect 25921 22811 26229 22820
rect 25261 22332 25569 22341
rect 25261 22330 25267 22332
rect 25323 22330 25347 22332
rect 25403 22330 25427 22332
rect 25483 22330 25507 22332
rect 25563 22330 25569 22332
rect 25323 22278 25325 22330
rect 25505 22278 25507 22330
rect 25261 22276 25267 22278
rect 25323 22276 25347 22278
rect 25403 22276 25427 22278
rect 25483 22276 25507 22278
rect 25563 22276 25569 22278
rect 25261 22267 25569 22276
rect 25921 21788 26229 21797
rect 25921 21786 25927 21788
rect 25983 21786 26007 21788
rect 26063 21786 26087 21788
rect 26143 21786 26167 21788
rect 26223 21786 26229 21788
rect 25983 21734 25985 21786
rect 26165 21734 26167 21786
rect 25921 21732 25927 21734
rect 25983 21732 26007 21734
rect 26063 21732 26087 21734
rect 26143 21732 26167 21734
rect 26223 21732 26229 21734
rect 25921 21723 26229 21732
rect 25261 21244 25569 21253
rect 25261 21242 25267 21244
rect 25323 21242 25347 21244
rect 25403 21242 25427 21244
rect 25483 21242 25507 21244
rect 25563 21242 25569 21244
rect 25323 21190 25325 21242
rect 25505 21190 25507 21242
rect 25261 21188 25267 21190
rect 25323 21188 25347 21190
rect 25403 21188 25427 21190
rect 25483 21188 25507 21190
rect 25563 21188 25569 21190
rect 25261 21179 25569 21188
rect 25921 20700 26229 20709
rect 25921 20698 25927 20700
rect 25983 20698 26007 20700
rect 26063 20698 26087 20700
rect 26143 20698 26167 20700
rect 26223 20698 26229 20700
rect 25983 20646 25985 20698
rect 26165 20646 26167 20698
rect 25921 20644 25927 20646
rect 25983 20644 26007 20646
rect 26063 20644 26087 20646
rect 26143 20644 26167 20646
rect 26223 20644 26229 20646
rect 25921 20635 26229 20644
rect 25261 20156 25569 20165
rect 25261 20154 25267 20156
rect 25323 20154 25347 20156
rect 25403 20154 25427 20156
rect 25483 20154 25507 20156
rect 25563 20154 25569 20156
rect 25323 20102 25325 20154
rect 25505 20102 25507 20154
rect 25261 20100 25267 20102
rect 25323 20100 25347 20102
rect 25403 20100 25427 20102
rect 25483 20100 25507 20102
rect 25563 20100 25569 20102
rect 25261 20091 25569 20100
rect 25921 19612 26229 19621
rect 25921 19610 25927 19612
rect 25983 19610 26007 19612
rect 26063 19610 26087 19612
rect 26143 19610 26167 19612
rect 26223 19610 26229 19612
rect 25983 19558 25985 19610
rect 26165 19558 26167 19610
rect 25921 19556 25927 19558
rect 25983 19556 26007 19558
rect 26063 19556 26087 19558
rect 26143 19556 26167 19558
rect 26223 19556 26229 19558
rect 25921 19547 26229 19556
rect 25261 19068 25569 19077
rect 25261 19066 25267 19068
rect 25323 19066 25347 19068
rect 25403 19066 25427 19068
rect 25483 19066 25507 19068
rect 25563 19066 25569 19068
rect 25323 19014 25325 19066
rect 25505 19014 25507 19066
rect 25261 19012 25267 19014
rect 25323 19012 25347 19014
rect 25403 19012 25427 19014
rect 25483 19012 25507 19014
rect 25563 19012 25569 19014
rect 25261 19003 25569 19012
rect 25921 18524 26229 18533
rect 25921 18522 25927 18524
rect 25983 18522 26007 18524
rect 26063 18522 26087 18524
rect 26143 18522 26167 18524
rect 26223 18522 26229 18524
rect 25983 18470 25985 18522
rect 26165 18470 26167 18522
rect 25921 18468 25927 18470
rect 25983 18468 26007 18470
rect 26063 18468 26087 18470
rect 26143 18468 26167 18470
rect 26223 18468 26229 18470
rect 25921 18459 26229 18468
rect 25261 17980 25569 17989
rect 25261 17978 25267 17980
rect 25323 17978 25347 17980
rect 25403 17978 25427 17980
rect 25483 17978 25507 17980
rect 25563 17978 25569 17980
rect 25323 17926 25325 17978
rect 25505 17926 25507 17978
rect 25261 17924 25267 17926
rect 25323 17924 25347 17926
rect 25403 17924 25427 17926
rect 25483 17924 25507 17926
rect 25563 17924 25569 17926
rect 25261 17915 25569 17924
rect 25921 17436 26229 17445
rect 25921 17434 25927 17436
rect 25983 17434 26007 17436
rect 26063 17434 26087 17436
rect 26143 17434 26167 17436
rect 26223 17434 26229 17436
rect 25983 17382 25985 17434
rect 26165 17382 26167 17434
rect 25921 17380 25927 17382
rect 25983 17380 26007 17382
rect 26063 17380 26087 17382
rect 26143 17380 26167 17382
rect 26223 17380 26229 17382
rect 25921 17371 26229 17380
rect 25261 16892 25569 16901
rect 25261 16890 25267 16892
rect 25323 16890 25347 16892
rect 25403 16890 25427 16892
rect 25483 16890 25507 16892
rect 25563 16890 25569 16892
rect 25323 16838 25325 16890
rect 25505 16838 25507 16890
rect 25261 16836 25267 16838
rect 25323 16836 25347 16838
rect 25403 16836 25427 16838
rect 25483 16836 25507 16838
rect 25563 16836 25569 16838
rect 25261 16827 25569 16836
rect 25921 16348 26229 16357
rect 25921 16346 25927 16348
rect 25983 16346 26007 16348
rect 26063 16346 26087 16348
rect 26143 16346 26167 16348
rect 26223 16346 26229 16348
rect 25983 16294 25985 16346
rect 26165 16294 26167 16346
rect 25921 16292 25927 16294
rect 25983 16292 26007 16294
rect 26063 16292 26087 16294
rect 26143 16292 26167 16294
rect 26223 16292 26229 16294
rect 25921 16283 26229 16292
rect 25261 15804 25569 15813
rect 25261 15802 25267 15804
rect 25323 15802 25347 15804
rect 25403 15802 25427 15804
rect 25483 15802 25507 15804
rect 25563 15802 25569 15804
rect 25323 15750 25325 15802
rect 25505 15750 25507 15802
rect 25261 15748 25267 15750
rect 25323 15748 25347 15750
rect 25403 15748 25427 15750
rect 25483 15748 25507 15750
rect 25563 15748 25569 15750
rect 25261 15739 25569 15748
rect 25921 15260 26229 15269
rect 25921 15258 25927 15260
rect 25983 15258 26007 15260
rect 26063 15258 26087 15260
rect 26143 15258 26167 15260
rect 26223 15258 26229 15260
rect 25983 15206 25985 15258
rect 26165 15206 26167 15258
rect 25921 15204 25927 15206
rect 25983 15204 26007 15206
rect 26063 15204 26087 15206
rect 26143 15204 26167 15206
rect 26223 15204 26229 15206
rect 25921 15195 26229 15204
rect 25261 14716 25569 14725
rect 25261 14714 25267 14716
rect 25323 14714 25347 14716
rect 25403 14714 25427 14716
rect 25483 14714 25507 14716
rect 25563 14714 25569 14716
rect 25323 14662 25325 14714
rect 25505 14662 25507 14714
rect 25261 14660 25267 14662
rect 25323 14660 25347 14662
rect 25403 14660 25427 14662
rect 25483 14660 25507 14662
rect 25563 14660 25569 14662
rect 25261 14651 25569 14660
rect 25921 14172 26229 14181
rect 25921 14170 25927 14172
rect 25983 14170 26007 14172
rect 26063 14170 26087 14172
rect 26143 14170 26167 14172
rect 26223 14170 26229 14172
rect 25983 14118 25985 14170
rect 26165 14118 26167 14170
rect 25921 14116 25927 14118
rect 25983 14116 26007 14118
rect 26063 14116 26087 14118
rect 26143 14116 26167 14118
rect 26223 14116 26229 14118
rect 25921 14107 26229 14116
rect 25261 13628 25569 13637
rect 25261 13626 25267 13628
rect 25323 13626 25347 13628
rect 25403 13626 25427 13628
rect 25483 13626 25507 13628
rect 25563 13626 25569 13628
rect 25323 13574 25325 13626
rect 25505 13574 25507 13626
rect 25261 13572 25267 13574
rect 25323 13572 25347 13574
rect 25403 13572 25427 13574
rect 25483 13572 25507 13574
rect 25563 13572 25569 13574
rect 25261 13563 25569 13572
rect 25921 13084 26229 13093
rect 25921 13082 25927 13084
rect 25983 13082 26007 13084
rect 26063 13082 26087 13084
rect 26143 13082 26167 13084
rect 26223 13082 26229 13084
rect 25983 13030 25985 13082
rect 26165 13030 26167 13082
rect 25921 13028 25927 13030
rect 25983 13028 26007 13030
rect 26063 13028 26087 13030
rect 26143 13028 26167 13030
rect 26223 13028 26229 13030
rect 25921 13019 26229 13028
rect 28276 12918 28304 25230
rect 28538 25191 28594 25200
rect 28264 12912 28316 12918
rect 28264 12854 28316 12860
rect 25261 12540 25569 12549
rect 25261 12538 25267 12540
rect 25323 12538 25347 12540
rect 25403 12538 25427 12540
rect 25483 12538 25507 12540
rect 25563 12538 25569 12540
rect 25323 12486 25325 12538
rect 25505 12486 25507 12538
rect 25261 12484 25267 12486
rect 25323 12484 25347 12486
rect 25403 12484 25427 12486
rect 25483 12484 25507 12486
rect 25563 12484 25569 12486
rect 25261 12475 25569 12484
rect 25921 11996 26229 12005
rect 25921 11994 25927 11996
rect 25983 11994 26007 11996
rect 26063 11994 26087 11996
rect 26143 11994 26167 11996
rect 26223 11994 26229 11996
rect 25983 11942 25985 11994
rect 26165 11942 26167 11994
rect 25921 11940 25927 11942
rect 25983 11940 26007 11942
rect 26063 11940 26087 11942
rect 26143 11940 26167 11942
rect 26223 11940 26229 11942
rect 25921 11931 26229 11940
rect 21732 11824 21784 11830
rect 21732 11766 21784 11772
rect 21640 11552 21692 11558
rect 21640 11494 21692 11500
rect 20996 11348 21048 11354
rect 20996 11290 21048 11296
rect 21456 11348 21508 11354
rect 21456 11290 21508 11296
rect 20720 11144 20772 11150
rect 20720 11086 20772 11092
rect 20732 10810 20760 11086
rect 20720 10804 20772 10810
rect 20720 10746 20772 10752
rect 20732 10130 20760 10746
rect 21272 10668 21324 10674
rect 21272 10610 21324 10616
rect 20812 10260 20864 10266
rect 20812 10202 20864 10208
rect 20720 10124 20772 10130
rect 20720 10066 20772 10072
rect 20260 9988 20312 9994
rect 20260 9930 20312 9936
rect 20168 9444 20220 9450
rect 20168 9386 20220 9392
rect 20272 9178 20300 9930
rect 20536 9920 20588 9926
rect 20536 9862 20588 9868
rect 20548 9518 20576 9862
rect 20824 9722 20852 10202
rect 21088 10056 21140 10062
rect 21088 9998 21140 10004
rect 21180 10056 21232 10062
rect 21180 9998 21232 10004
rect 20904 9920 20956 9926
rect 20904 9862 20956 9868
rect 20812 9716 20864 9722
rect 20812 9658 20864 9664
rect 20916 9586 20944 9862
rect 20904 9580 20956 9586
rect 20904 9522 20956 9528
rect 20996 9580 21048 9586
rect 20996 9522 21048 9528
rect 20536 9512 20588 9518
rect 20536 9454 20588 9460
rect 21008 9382 21036 9522
rect 21100 9450 21128 9998
rect 21088 9444 21140 9450
rect 21088 9386 21140 9392
rect 20812 9376 20864 9382
rect 20812 9318 20864 9324
rect 20996 9376 21048 9382
rect 20996 9318 21048 9324
rect 20260 9172 20312 9178
rect 20260 9114 20312 9120
rect 20720 9172 20772 9178
rect 20720 9114 20772 9120
rect 20352 8832 20404 8838
rect 20352 8774 20404 8780
rect 20536 8832 20588 8838
rect 20536 8774 20588 8780
rect 20364 8634 20392 8774
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 20260 8492 20312 8498
rect 20260 8434 20312 8440
rect 20168 8424 20220 8430
rect 20168 8366 20220 8372
rect 20076 7880 20128 7886
rect 20076 7822 20128 7828
rect 20180 7818 20208 8366
rect 20272 8090 20300 8434
rect 20548 8430 20576 8774
rect 20536 8424 20588 8430
rect 20536 8366 20588 8372
rect 20260 8084 20312 8090
rect 20260 8026 20312 8032
rect 20732 8022 20760 9114
rect 20824 9110 20852 9318
rect 20812 9104 20864 9110
rect 20812 9046 20864 9052
rect 20824 8634 20852 9046
rect 20904 9036 20956 9042
rect 20904 8978 20956 8984
rect 20812 8628 20864 8634
rect 20812 8570 20864 8576
rect 20720 8016 20772 8022
rect 20720 7958 20772 7964
rect 20812 8016 20864 8022
rect 20812 7958 20864 7964
rect 20168 7812 20220 7818
rect 20168 7754 20220 7760
rect 20444 7812 20496 7818
rect 20444 7754 20496 7760
rect 20456 7478 20484 7754
rect 20732 7750 20760 7958
rect 20720 7744 20772 7750
rect 20720 7686 20772 7692
rect 20732 7546 20760 7686
rect 20720 7540 20772 7546
rect 20720 7482 20772 7488
rect 19708 7472 19760 7478
rect 19708 7414 19760 7420
rect 20444 7472 20496 7478
rect 20444 7414 20496 7420
rect 18236 6656 18288 6662
rect 18236 6598 18288 6604
rect 18248 6390 18276 6598
rect 18236 6384 18288 6390
rect 18236 6326 18288 6332
rect 18064 5902 18184 5930
rect 17868 5704 17920 5710
rect 17868 5646 17920 5652
rect 17960 5568 18012 5574
rect 17960 5510 18012 5516
rect 17408 4820 17460 4826
rect 17408 4762 17460 4768
rect 17972 4622 18000 5510
rect 18052 5024 18104 5030
rect 18052 4966 18104 4972
rect 17960 4616 18012 4622
rect 17960 4558 18012 4564
rect 17960 4480 18012 4486
rect 17960 4422 18012 4428
rect 17408 3936 17460 3942
rect 17408 3878 17460 3884
rect 17420 3194 17448 3878
rect 17972 3534 18000 4422
rect 18064 4078 18092 4966
rect 18052 4072 18104 4078
rect 18052 4014 18104 4020
rect 17868 3528 17920 3534
rect 17868 3470 17920 3476
rect 17960 3528 18012 3534
rect 17960 3470 18012 3476
rect 17408 3188 17460 3194
rect 17408 3130 17460 3136
rect 17880 3058 17908 3470
rect 17868 3052 17920 3058
rect 17868 2994 17920 3000
rect 17144 2746 17264 2774
rect 13544 2508 13596 2514
rect 13544 2450 13596 2456
rect 20 2440 72 2446
rect 20 2382 72 2388
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 32 800 60 2382
rect 5083 2204 5391 2213
rect 5083 2202 5089 2204
rect 5145 2202 5169 2204
rect 5225 2202 5249 2204
rect 5305 2202 5329 2204
rect 5385 2202 5391 2204
rect 5145 2150 5147 2202
rect 5327 2150 5329 2202
rect 5083 2148 5089 2150
rect 5145 2148 5169 2150
rect 5225 2148 5249 2150
rect 5305 2148 5329 2150
rect 5385 2148 5391 2150
rect 5083 2139 5391 2148
rect 9140 1306 9168 2382
rect 17144 2378 17172 2746
rect 18156 2650 18184 5902
rect 18248 5352 18276 6326
rect 18315 6012 18623 6021
rect 18315 6010 18321 6012
rect 18377 6010 18401 6012
rect 18457 6010 18481 6012
rect 18537 6010 18561 6012
rect 18617 6010 18623 6012
rect 18377 5958 18379 6010
rect 18559 5958 18561 6010
rect 18315 5956 18321 5958
rect 18377 5956 18401 5958
rect 18457 5956 18481 5958
rect 18537 5956 18561 5958
rect 18617 5956 18623 5958
rect 18315 5947 18623 5956
rect 18248 5324 18368 5352
rect 18236 5228 18288 5234
rect 18236 5170 18288 5176
rect 18248 4826 18276 5170
rect 18340 5166 18368 5324
rect 18328 5160 18380 5166
rect 18328 5102 18380 5108
rect 18315 4924 18623 4933
rect 18315 4922 18321 4924
rect 18377 4922 18401 4924
rect 18457 4922 18481 4924
rect 18537 4922 18561 4924
rect 18617 4922 18623 4924
rect 18377 4870 18379 4922
rect 18559 4870 18561 4922
rect 18315 4868 18321 4870
rect 18377 4868 18401 4870
rect 18457 4868 18481 4870
rect 18537 4868 18561 4870
rect 18617 4868 18623 4870
rect 18315 4859 18623 4868
rect 18236 4820 18288 4826
rect 18236 4762 18288 4768
rect 18708 4078 18736 6734
rect 18800 6718 18920 6746
rect 18788 6656 18840 6662
rect 18788 6598 18840 6604
rect 18800 5302 18828 6598
rect 18788 5296 18840 5302
rect 18788 5238 18840 5244
rect 18892 4758 18920 6718
rect 18975 6556 19283 6565
rect 18975 6554 18981 6556
rect 19037 6554 19061 6556
rect 19117 6554 19141 6556
rect 19197 6554 19221 6556
rect 19277 6554 19283 6556
rect 19037 6502 19039 6554
rect 19219 6502 19221 6554
rect 18975 6500 18981 6502
rect 19037 6500 19061 6502
rect 19117 6500 19141 6502
rect 19197 6500 19221 6502
rect 19277 6500 19283 6502
rect 18975 6491 19283 6500
rect 19720 6390 19748 7414
rect 19708 6384 19760 6390
rect 19708 6326 19760 6332
rect 20732 6322 20760 7482
rect 20824 7313 20852 7958
rect 20916 7886 20944 8978
rect 20996 8968 21048 8974
rect 20996 8910 21048 8916
rect 21008 7954 21036 8910
rect 21100 8498 21128 9386
rect 21192 9382 21220 9998
rect 21180 9376 21232 9382
rect 21180 9318 21232 9324
rect 21088 8492 21140 8498
rect 21088 8434 21140 8440
rect 21192 8430 21220 9318
rect 21284 9178 21312 10610
rect 21364 10192 21416 10198
rect 21364 10134 21416 10140
rect 21376 9654 21404 10134
rect 21364 9648 21416 9654
rect 21364 9590 21416 9596
rect 21272 9172 21324 9178
rect 21272 9114 21324 9120
rect 21376 8974 21404 9590
rect 21468 8974 21496 11290
rect 21548 10464 21600 10470
rect 21548 10406 21600 10412
rect 21560 9994 21588 10406
rect 21652 10130 21680 11494
rect 21640 10124 21692 10130
rect 21640 10066 21692 10072
rect 21548 9988 21600 9994
rect 21600 9948 21680 9976
rect 21548 9930 21600 9936
rect 21652 9586 21680 9948
rect 21640 9580 21692 9586
rect 21640 9522 21692 9528
rect 21364 8968 21416 8974
rect 21364 8910 21416 8916
rect 21456 8968 21508 8974
rect 21456 8910 21508 8916
rect 21456 8832 21508 8838
rect 21456 8774 21508 8780
rect 21548 8832 21600 8838
rect 21548 8774 21600 8780
rect 21468 8498 21496 8774
rect 21560 8634 21588 8774
rect 21548 8628 21600 8634
rect 21548 8570 21600 8576
rect 21652 8498 21680 9522
rect 21456 8492 21508 8498
rect 21456 8434 21508 8440
rect 21640 8492 21692 8498
rect 21640 8434 21692 8440
rect 21180 8424 21232 8430
rect 21180 8366 21232 8372
rect 21192 8090 21220 8366
rect 21180 8084 21232 8090
rect 21180 8026 21232 8032
rect 20996 7948 21048 7954
rect 20996 7890 21048 7896
rect 20904 7880 20956 7886
rect 20904 7822 20956 7828
rect 20810 7304 20866 7313
rect 20916 7274 20944 7822
rect 21008 7546 21036 7890
rect 20996 7540 21048 7546
rect 20996 7482 21048 7488
rect 21192 7410 21220 8026
rect 21468 7478 21496 8434
rect 21456 7472 21508 7478
rect 21456 7414 21508 7420
rect 21180 7404 21232 7410
rect 21180 7346 21232 7352
rect 21640 7404 21692 7410
rect 21640 7346 21692 7352
rect 20810 7239 20866 7248
rect 20904 7268 20956 7274
rect 20536 6316 20588 6322
rect 20536 6258 20588 6264
rect 20720 6316 20772 6322
rect 20720 6258 20772 6264
rect 19340 6248 19392 6254
rect 19340 6190 19392 6196
rect 19352 5846 19380 6190
rect 19800 6112 19852 6118
rect 19800 6054 19852 6060
rect 20168 6112 20220 6118
rect 20168 6054 20220 6060
rect 19340 5840 19392 5846
rect 19340 5782 19392 5788
rect 18975 5468 19283 5477
rect 18975 5466 18981 5468
rect 19037 5466 19061 5468
rect 19117 5466 19141 5468
rect 19197 5466 19221 5468
rect 19277 5466 19283 5468
rect 19037 5414 19039 5466
rect 19219 5414 19221 5466
rect 18975 5412 18981 5414
rect 19037 5412 19061 5414
rect 19117 5412 19141 5414
rect 19197 5412 19221 5414
rect 19277 5412 19283 5414
rect 18975 5403 19283 5412
rect 18972 5092 19024 5098
rect 18972 5034 19024 5040
rect 18880 4752 18932 4758
rect 18880 4694 18932 4700
rect 18788 4616 18840 4622
rect 18788 4558 18840 4564
rect 18696 4072 18748 4078
rect 18696 4014 18748 4020
rect 18315 3836 18623 3845
rect 18315 3834 18321 3836
rect 18377 3834 18401 3836
rect 18457 3834 18481 3836
rect 18537 3834 18561 3836
rect 18617 3834 18623 3836
rect 18377 3782 18379 3834
rect 18559 3782 18561 3834
rect 18315 3780 18321 3782
rect 18377 3780 18401 3782
rect 18457 3780 18481 3782
rect 18537 3780 18561 3782
rect 18617 3780 18623 3782
rect 18315 3771 18623 3780
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 18616 3126 18644 3470
rect 18604 3120 18656 3126
rect 18604 3062 18656 3068
rect 18315 2748 18623 2757
rect 18315 2746 18321 2748
rect 18377 2746 18401 2748
rect 18457 2746 18481 2748
rect 18537 2746 18561 2748
rect 18617 2746 18623 2748
rect 18377 2694 18379 2746
rect 18559 2694 18561 2746
rect 18315 2692 18321 2694
rect 18377 2692 18401 2694
rect 18457 2692 18481 2694
rect 18537 2692 18561 2694
rect 18617 2692 18623 2694
rect 18315 2683 18623 2692
rect 18144 2644 18196 2650
rect 18144 2586 18196 2592
rect 18052 2440 18104 2446
rect 18052 2382 18104 2388
rect 17132 2372 17184 2378
rect 17132 2314 17184 2320
rect 12029 2204 12337 2213
rect 12029 2202 12035 2204
rect 12091 2202 12115 2204
rect 12171 2202 12195 2204
rect 12251 2202 12275 2204
rect 12331 2202 12337 2204
rect 12091 2150 12093 2202
rect 12273 2150 12275 2202
rect 12029 2148 12035 2150
rect 12091 2148 12115 2150
rect 12171 2148 12195 2150
rect 12251 2148 12275 2150
rect 12331 2148 12337 2150
rect 12029 2139 12337 2148
rect 9048 1278 9168 1306
rect 9048 800 9076 1278
rect 18064 800 18092 2382
rect 18800 2310 18828 4558
rect 18892 3398 18920 4694
rect 18984 4622 19012 5034
rect 19352 5030 19380 5782
rect 19812 5778 19840 6054
rect 19800 5772 19852 5778
rect 19800 5714 19852 5720
rect 19812 5658 19840 5714
rect 20180 5710 20208 6054
rect 20548 5914 20576 6258
rect 20536 5908 20588 5914
rect 20536 5850 20588 5856
rect 19720 5630 19840 5658
rect 20076 5704 20128 5710
rect 20076 5646 20128 5652
rect 20168 5704 20220 5710
rect 20168 5646 20220 5652
rect 19432 5228 19484 5234
rect 19432 5170 19484 5176
rect 19340 5024 19392 5030
rect 19340 4966 19392 4972
rect 19340 4820 19392 4826
rect 19340 4762 19392 4768
rect 18972 4616 19024 4622
rect 18972 4558 19024 4564
rect 18975 4380 19283 4389
rect 18975 4378 18981 4380
rect 19037 4378 19061 4380
rect 19117 4378 19141 4380
rect 19197 4378 19221 4380
rect 19277 4378 19283 4380
rect 19037 4326 19039 4378
rect 19219 4326 19221 4378
rect 18975 4324 18981 4326
rect 19037 4324 19061 4326
rect 19117 4324 19141 4326
rect 19197 4324 19221 4326
rect 19277 4324 19283 4326
rect 18975 4315 19283 4324
rect 18970 4176 19026 4185
rect 19352 4146 19380 4762
rect 19444 4146 19472 5170
rect 19720 5030 19748 5630
rect 19800 5568 19852 5574
rect 19800 5510 19852 5516
rect 19708 5024 19760 5030
rect 19708 4966 19760 4972
rect 19524 4548 19576 4554
rect 19524 4490 19576 4496
rect 19616 4548 19668 4554
rect 19616 4490 19668 4496
rect 19536 4282 19564 4490
rect 19524 4276 19576 4282
rect 19524 4218 19576 4224
rect 18970 4111 18972 4120
rect 19024 4111 19026 4120
rect 19340 4140 19392 4146
rect 18972 4082 19024 4088
rect 19340 4082 19392 4088
rect 19432 4140 19484 4146
rect 19432 4082 19484 4088
rect 19444 3738 19472 4082
rect 19628 3754 19656 4490
rect 19812 4486 19840 5510
rect 20088 5250 20116 5646
rect 20088 5234 20300 5250
rect 19892 5228 19944 5234
rect 20088 5228 20312 5234
rect 20088 5222 20260 5228
rect 19892 5170 19944 5176
rect 20260 5170 20312 5176
rect 19800 4480 19852 4486
rect 19800 4422 19852 4428
rect 19812 4078 19840 4422
rect 19800 4072 19852 4078
rect 19800 4014 19852 4020
rect 19708 3936 19760 3942
rect 19708 3878 19760 3884
rect 19432 3732 19484 3738
rect 19432 3674 19484 3680
rect 19536 3726 19656 3754
rect 18880 3392 18932 3398
rect 18880 3334 18932 3340
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 18975 3292 19283 3301
rect 18975 3290 18981 3292
rect 19037 3290 19061 3292
rect 19117 3290 19141 3292
rect 19197 3290 19221 3292
rect 19277 3290 19283 3292
rect 19037 3238 19039 3290
rect 19219 3238 19221 3290
rect 18975 3236 18981 3238
rect 19037 3236 19061 3238
rect 19117 3236 19141 3238
rect 19197 3236 19221 3238
rect 19277 3236 19283 3238
rect 18975 3227 19283 3236
rect 19352 2514 19380 3334
rect 19536 3194 19564 3726
rect 19616 3596 19668 3602
rect 19616 3538 19668 3544
rect 19628 3194 19656 3538
rect 19524 3188 19576 3194
rect 19524 3130 19576 3136
rect 19616 3188 19668 3194
rect 19616 3130 19668 3136
rect 19720 2774 19748 3878
rect 19812 3194 19840 4014
rect 19904 3602 19932 5170
rect 20272 3942 20300 5170
rect 20352 5024 20404 5030
rect 20352 4966 20404 4972
rect 20364 4282 20392 4966
rect 20352 4276 20404 4282
rect 20352 4218 20404 4224
rect 20260 3936 20312 3942
rect 20260 3878 20312 3884
rect 19892 3596 19944 3602
rect 19892 3538 19944 3544
rect 20272 3534 20300 3878
rect 20824 3534 20852 7239
rect 20904 7210 20956 7216
rect 21180 7200 21232 7206
rect 21180 7142 21232 7148
rect 21192 6322 21220 7142
rect 21180 6316 21232 6322
rect 21180 6258 21232 6264
rect 21652 5234 21680 7346
rect 21744 6712 21772 11766
rect 25261 11452 25569 11461
rect 25261 11450 25267 11452
rect 25323 11450 25347 11452
rect 25403 11450 25427 11452
rect 25483 11450 25507 11452
rect 25563 11450 25569 11452
rect 25323 11398 25325 11450
rect 25505 11398 25507 11450
rect 25261 11396 25267 11398
rect 25323 11396 25347 11398
rect 25403 11396 25427 11398
rect 25483 11396 25507 11398
rect 25563 11396 25569 11398
rect 25261 11387 25569 11396
rect 22008 11076 22060 11082
rect 22008 11018 22060 11024
rect 22468 11076 22520 11082
rect 22468 11018 22520 11024
rect 21824 10668 21876 10674
rect 21824 10610 21876 10616
rect 21836 10062 21864 10610
rect 21916 10532 21968 10538
rect 21916 10474 21968 10480
rect 21824 10056 21876 10062
rect 21824 9998 21876 10004
rect 21928 9722 21956 10474
rect 22020 10266 22048 11018
rect 22480 10810 22508 11018
rect 22560 11008 22612 11014
rect 22560 10950 22612 10956
rect 22468 10804 22520 10810
rect 22468 10746 22520 10752
rect 22284 10668 22336 10674
rect 22284 10610 22336 10616
rect 22008 10260 22060 10266
rect 22008 10202 22060 10208
rect 22008 10056 22060 10062
rect 22008 9998 22060 10004
rect 21916 9716 21968 9722
rect 21836 9676 21916 9704
rect 21836 8974 21864 9676
rect 21916 9658 21968 9664
rect 22020 9654 22048 9998
rect 22296 9722 22324 10610
rect 22572 10606 22600 10950
rect 25921 10908 26229 10917
rect 25921 10906 25927 10908
rect 25983 10906 26007 10908
rect 26063 10906 26087 10908
rect 26143 10906 26167 10908
rect 26223 10906 26229 10908
rect 25983 10854 25985 10906
rect 26165 10854 26167 10906
rect 25921 10852 25927 10854
rect 25983 10852 26007 10854
rect 26063 10852 26087 10854
rect 26143 10852 26167 10854
rect 26223 10852 26229 10854
rect 25921 10843 26229 10852
rect 23940 10804 23992 10810
rect 23940 10746 23992 10752
rect 22560 10600 22612 10606
rect 22560 10542 22612 10548
rect 22572 10130 22600 10542
rect 22560 10124 22612 10130
rect 22560 10066 22612 10072
rect 23204 10124 23256 10130
rect 23204 10066 23256 10072
rect 22468 9988 22520 9994
rect 22468 9930 22520 9936
rect 22480 9722 22508 9930
rect 22560 9920 22612 9926
rect 22560 9862 22612 9868
rect 22284 9716 22336 9722
rect 22284 9658 22336 9664
rect 22468 9716 22520 9722
rect 22468 9658 22520 9664
rect 22008 9648 22060 9654
rect 22008 9590 22060 9596
rect 22284 9376 22336 9382
rect 22284 9318 22336 9324
rect 22296 9178 22324 9318
rect 22284 9172 22336 9178
rect 22284 9114 22336 9120
rect 22008 9104 22060 9110
rect 22008 9046 22060 9052
rect 21824 8968 21876 8974
rect 21824 8910 21876 8916
rect 22020 8634 22048 9046
rect 22468 8832 22520 8838
rect 22468 8774 22520 8780
rect 22008 8628 22060 8634
rect 22008 8570 22060 8576
rect 21822 8256 21878 8265
rect 21822 8191 21878 8200
rect 21836 7886 21864 8191
rect 22480 8022 22508 8774
rect 22572 8498 22600 9862
rect 22652 9512 22704 9518
rect 22652 9454 22704 9460
rect 22664 8974 22692 9454
rect 22652 8968 22704 8974
rect 22652 8910 22704 8916
rect 22836 8900 22888 8906
rect 22836 8842 22888 8848
rect 22652 8832 22704 8838
rect 22652 8774 22704 8780
rect 22664 8634 22692 8774
rect 22652 8628 22704 8634
rect 22652 8570 22704 8576
rect 22560 8492 22612 8498
rect 22560 8434 22612 8440
rect 22468 8016 22520 8022
rect 22468 7958 22520 7964
rect 21824 7880 21876 7886
rect 21824 7822 21876 7828
rect 22480 7546 22508 7958
rect 22560 7744 22612 7750
rect 22560 7686 22612 7692
rect 22468 7540 22520 7546
rect 22468 7482 22520 7488
rect 21916 7404 21968 7410
rect 21916 7346 21968 7352
rect 22192 7404 22244 7410
rect 22192 7346 22244 7352
rect 21928 7313 21956 7346
rect 21914 7304 21970 7313
rect 21914 7239 21970 7248
rect 21824 6724 21876 6730
rect 21744 6684 21824 6712
rect 21744 5710 21772 6684
rect 21824 6666 21876 6672
rect 21732 5704 21784 5710
rect 21732 5646 21784 5652
rect 20996 5228 21048 5234
rect 20996 5170 21048 5176
rect 21640 5228 21692 5234
rect 21640 5170 21692 5176
rect 21008 4826 21036 5170
rect 20996 4820 21048 4826
rect 20996 4762 21048 4768
rect 21272 4616 21324 4622
rect 21272 4558 21324 4564
rect 21456 4616 21508 4622
rect 21456 4558 21508 4564
rect 20260 3528 20312 3534
rect 20260 3470 20312 3476
rect 20812 3528 20864 3534
rect 20812 3470 20864 3476
rect 20904 3460 20956 3466
rect 20904 3402 20956 3408
rect 20720 3392 20772 3398
rect 20720 3334 20772 3340
rect 19800 3188 19852 3194
rect 19800 3130 19852 3136
rect 19984 2984 20036 2990
rect 19984 2926 20036 2932
rect 19628 2746 19748 2774
rect 19340 2508 19392 2514
rect 19340 2450 19392 2456
rect 19628 2446 19656 2746
rect 19996 2650 20024 2926
rect 19984 2644 20036 2650
rect 19984 2586 20036 2592
rect 20732 2446 20760 3334
rect 20916 2446 20944 3402
rect 21180 2984 21232 2990
rect 21180 2926 21232 2932
rect 21192 2650 21220 2926
rect 21284 2650 21312 4558
rect 21468 3738 21496 4558
rect 21548 4480 21600 4486
rect 21548 4422 21600 4428
rect 21560 4282 21588 4422
rect 21548 4276 21600 4282
rect 21548 4218 21600 4224
rect 21744 4214 21772 5646
rect 21928 5370 21956 7239
rect 22204 6798 22232 7346
rect 22572 7342 22600 7686
rect 22376 7336 22428 7342
rect 22376 7278 22428 7284
rect 22560 7336 22612 7342
rect 22560 7278 22612 7284
rect 22388 7188 22416 7278
rect 22560 7200 22612 7206
rect 22388 7160 22560 7188
rect 22560 7142 22612 7148
rect 22192 6792 22244 6798
rect 22664 6746 22692 8570
rect 22848 8090 22876 8842
rect 23216 8430 23244 10066
rect 23388 9444 23440 9450
rect 23388 9386 23440 9392
rect 23400 8974 23428 9386
rect 23388 8968 23440 8974
rect 23388 8910 23440 8916
rect 23400 8634 23428 8910
rect 23480 8832 23532 8838
rect 23480 8774 23532 8780
rect 23756 8832 23808 8838
rect 23756 8774 23808 8780
rect 23388 8628 23440 8634
rect 23388 8570 23440 8576
rect 23492 8566 23520 8774
rect 23768 8634 23796 8774
rect 23756 8628 23808 8634
rect 23756 8570 23808 8576
rect 23480 8560 23532 8566
rect 23480 8502 23532 8508
rect 23204 8424 23256 8430
rect 23204 8366 23256 8372
rect 22836 8084 22888 8090
rect 22836 8026 22888 8032
rect 23216 7750 23244 8366
rect 23492 8090 23520 8502
rect 23952 8090 23980 10746
rect 24032 10668 24084 10674
rect 24032 10610 24084 10616
rect 24044 9994 24072 10610
rect 24308 10464 24360 10470
rect 24308 10406 24360 10412
rect 24320 9994 24348 10406
rect 25261 10364 25569 10373
rect 25261 10362 25267 10364
rect 25323 10362 25347 10364
rect 25403 10362 25427 10364
rect 25483 10362 25507 10364
rect 25563 10362 25569 10364
rect 25323 10310 25325 10362
rect 25505 10310 25507 10362
rect 25261 10308 25267 10310
rect 25323 10308 25347 10310
rect 25403 10308 25427 10310
rect 25483 10308 25507 10310
rect 25563 10308 25569 10310
rect 25261 10299 25569 10308
rect 24032 9988 24084 9994
rect 24032 9930 24084 9936
rect 24308 9988 24360 9994
rect 24308 9930 24360 9936
rect 24044 8566 24072 9930
rect 24124 9512 24176 9518
rect 24124 9454 24176 9460
rect 24136 8838 24164 9454
rect 24124 8832 24176 8838
rect 24124 8774 24176 8780
rect 24032 8560 24084 8566
rect 24032 8502 24084 8508
rect 23480 8084 23532 8090
rect 23480 8026 23532 8032
rect 23940 8084 23992 8090
rect 23940 8026 23992 8032
rect 23952 7970 23980 8026
rect 23952 7954 24072 7970
rect 24136 7954 24164 8774
rect 24216 8288 24268 8294
rect 24216 8230 24268 8236
rect 23952 7948 24084 7954
rect 23952 7942 24032 7948
rect 24032 7890 24084 7896
rect 24124 7948 24176 7954
rect 24124 7890 24176 7896
rect 24228 7818 24256 8230
rect 24216 7812 24268 7818
rect 24216 7754 24268 7760
rect 24320 7750 24348 9930
rect 25921 9820 26229 9829
rect 25921 9818 25927 9820
rect 25983 9818 26007 9820
rect 26063 9818 26087 9820
rect 26143 9818 26167 9820
rect 26223 9818 26229 9820
rect 25983 9766 25985 9818
rect 26165 9766 26167 9818
rect 25921 9764 25927 9766
rect 25983 9764 26007 9766
rect 26063 9764 26087 9766
rect 26143 9764 26167 9766
rect 26223 9764 26229 9766
rect 25921 9755 26229 9764
rect 25261 9276 25569 9285
rect 25261 9274 25267 9276
rect 25323 9274 25347 9276
rect 25403 9274 25427 9276
rect 25483 9274 25507 9276
rect 25563 9274 25569 9276
rect 25323 9222 25325 9274
rect 25505 9222 25507 9274
rect 25261 9220 25267 9222
rect 25323 9220 25347 9222
rect 25403 9220 25427 9222
rect 25483 9220 25507 9222
rect 25563 9220 25569 9222
rect 25261 9211 25569 9220
rect 24768 8968 24820 8974
rect 24768 8910 24820 8916
rect 24780 8294 24808 8910
rect 25921 8732 26229 8741
rect 25921 8730 25927 8732
rect 25983 8730 26007 8732
rect 26063 8730 26087 8732
rect 26143 8730 26167 8732
rect 26223 8730 26229 8732
rect 25983 8678 25985 8730
rect 26165 8678 26167 8730
rect 25921 8676 25927 8678
rect 25983 8676 26007 8678
rect 26063 8676 26087 8678
rect 26143 8676 26167 8678
rect 26223 8676 26229 8678
rect 25921 8667 26229 8676
rect 24768 8288 24820 8294
rect 24768 8230 24820 8236
rect 24780 8090 24808 8230
rect 25261 8188 25569 8197
rect 25261 8186 25267 8188
rect 25323 8186 25347 8188
rect 25403 8186 25427 8188
rect 25483 8186 25507 8188
rect 25563 8186 25569 8188
rect 25323 8134 25325 8186
rect 25505 8134 25507 8186
rect 25261 8132 25267 8134
rect 25323 8132 25347 8134
rect 25403 8132 25427 8134
rect 25483 8132 25507 8134
rect 25563 8132 25569 8134
rect 25261 8123 25569 8132
rect 24768 8084 24820 8090
rect 24768 8026 24820 8032
rect 28264 7812 28316 7818
rect 28264 7754 28316 7760
rect 23204 7744 23256 7750
rect 23204 7686 23256 7692
rect 24308 7744 24360 7750
rect 24308 7686 24360 7692
rect 24860 7744 24912 7750
rect 24860 7686 24912 7692
rect 25044 7744 25096 7750
rect 25044 7686 25096 7692
rect 23216 7342 23244 7686
rect 24872 7392 24900 7686
rect 24780 7364 24900 7392
rect 22744 7336 22796 7342
rect 22744 7278 22796 7284
rect 22836 7336 22888 7342
rect 23020 7336 23072 7342
rect 22940 7313 23020 7324
rect 22836 7278 22888 7284
rect 22926 7304 23020 7313
rect 22192 6734 22244 6740
rect 22204 6458 22232 6734
rect 22376 6724 22428 6730
rect 22376 6666 22428 6672
rect 22572 6718 22692 6746
rect 22192 6452 22244 6458
rect 22192 6394 22244 6400
rect 22192 6316 22244 6322
rect 22192 6258 22244 6264
rect 22204 5642 22232 6258
rect 22388 6186 22416 6666
rect 22376 6180 22428 6186
rect 22376 6122 22428 6128
rect 22388 5710 22416 6122
rect 22572 6118 22600 6718
rect 22652 6656 22704 6662
rect 22652 6598 22704 6604
rect 22664 6458 22692 6598
rect 22652 6452 22704 6458
rect 22652 6394 22704 6400
rect 22560 6112 22612 6118
rect 22560 6054 22612 6060
rect 22376 5704 22428 5710
rect 22376 5646 22428 5652
rect 22100 5636 22152 5642
rect 22100 5578 22152 5584
rect 22192 5636 22244 5642
rect 22192 5578 22244 5584
rect 22284 5636 22336 5642
rect 22284 5578 22336 5584
rect 22112 5370 22140 5578
rect 22204 5370 22232 5578
rect 21916 5364 21968 5370
rect 21916 5306 21968 5312
rect 22100 5364 22152 5370
rect 22100 5306 22152 5312
rect 22192 5364 22244 5370
rect 22192 5306 22244 5312
rect 22296 5302 22324 5578
rect 22284 5296 22336 5302
rect 22284 5238 22336 5244
rect 22284 5024 22336 5030
rect 22284 4966 22336 4972
rect 22296 4826 22324 4966
rect 22284 4820 22336 4826
rect 22284 4762 22336 4768
rect 21916 4480 21968 4486
rect 21916 4422 21968 4428
rect 21928 4282 21956 4422
rect 21916 4276 21968 4282
rect 21916 4218 21968 4224
rect 21732 4208 21784 4214
rect 21732 4150 21784 4156
rect 22192 4208 22244 4214
rect 22388 4196 22416 5646
rect 22468 5636 22520 5642
rect 22468 5578 22520 5584
rect 22480 5098 22508 5578
rect 22468 5092 22520 5098
rect 22468 5034 22520 5040
rect 22480 4282 22508 5034
rect 22468 4276 22520 4282
rect 22468 4218 22520 4224
rect 22244 4168 22416 4196
rect 22192 4150 22244 4156
rect 21456 3732 21508 3738
rect 21456 3674 21508 3680
rect 21468 2922 21496 3674
rect 21744 3126 21772 4150
rect 22204 3738 22232 4150
rect 22192 3732 22244 3738
rect 22192 3674 22244 3680
rect 22572 3466 22600 6054
rect 22756 5914 22784 7278
rect 22848 6390 22876 7278
rect 22982 7296 23020 7304
rect 23020 7278 23072 7284
rect 23204 7336 23256 7342
rect 23204 7278 23256 7284
rect 23664 7336 23716 7342
rect 23664 7278 23716 7284
rect 22926 7239 22982 7248
rect 23216 6866 23244 7278
rect 23676 7002 23704 7278
rect 23664 6996 23716 7002
rect 23664 6938 23716 6944
rect 23572 6928 23624 6934
rect 23572 6870 23624 6876
rect 23204 6860 23256 6866
rect 23204 6802 23256 6808
rect 23480 6792 23532 6798
rect 23480 6734 23532 6740
rect 23296 6656 23348 6662
rect 23296 6598 23348 6604
rect 23204 6452 23256 6458
rect 23204 6394 23256 6400
rect 22836 6384 22888 6390
rect 22836 6326 22888 6332
rect 23020 6316 23072 6322
rect 23020 6258 23072 6264
rect 22744 5908 22796 5914
rect 22744 5850 22796 5856
rect 23032 5778 23060 6258
rect 23020 5772 23072 5778
rect 23020 5714 23072 5720
rect 23216 5370 23244 6394
rect 23308 6322 23336 6598
rect 23296 6316 23348 6322
rect 23296 6258 23348 6264
rect 23492 6254 23520 6734
rect 23584 6458 23612 6870
rect 23756 6792 23808 6798
rect 23756 6734 23808 6740
rect 23768 6458 23796 6734
rect 23572 6452 23624 6458
rect 23572 6394 23624 6400
rect 23756 6452 23808 6458
rect 23756 6394 23808 6400
rect 24780 6390 24808 7364
rect 24860 7268 24912 7274
rect 24860 7210 24912 7216
rect 24872 6474 24900 7210
rect 24952 7200 25004 7206
rect 24952 7142 25004 7148
rect 24964 6866 24992 7142
rect 25056 7002 25084 7686
rect 25921 7644 26229 7653
rect 25921 7642 25927 7644
rect 25983 7642 26007 7644
rect 26063 7642 26087 7644
rect 26143 7642 26167 7644
rect 26223 7642 26229 7644
rect 25983 7590 25985 7642
rect 26165 7590 26167 7642
rect 25921 7588 25927 7590
rect 25983 7588 26007 7590
rect 26063 7588 26087 7590
rect 26143 7588 26167 7590
rect 26223 7588 26229 7590
rect 25921 7579 26229 7588
rect 25261 7100 25569 7109
rect 25261 7098 25267 7100
rect 25323 7098 25347 7100
rect 25403 7098 25427 7100
rect 25483 7098 25507 7100
rect 25563 7098 25569 7100
rect 25323 7046 25325 7098
rect 25505 7046 25507 7098
rect 25261 7044 25267 7046
rect 25323 7044 25347 7046
rect 25403 7044 25427 7046
rect 25483 7044 25507 7046
rect 25563 7044 25569 7046
rect 25261 7035 25569 7044
rect 25044 6996 25096 7002
rect 25044 6938 25096 6944
rect 25596 6996 25648 7002
rect 25596 6938 25648 6944
rect 24952 6860 25004 6866
rect 24952 6802 25004 6808
rect 25056 6662 25084 6938
rect 25044 6656 25096 6662
rect 25044 6598 25096 6604
rect 25136 6656 25188 6662
rect 25136 6598 25188 6604
rect 25504 6656 25556 6662
rect 25504 6598 25556 6604
rect 24872 6446 24992 6474
rect 24964 6390 24992 6446
rect 24768 6384 24820 6390
rect 24768 6326 24820 6332
rect 24952 6384 25004 6390
rect 24952 6326 25004 6332
rect 23848 6316 23900 6322
rect 23848 6258 23900 6264
rect 24032 6316 24084 6322
rect 24032 6258 24084 6264
rect 23480 6248 23532 6254
rect 23480 6190 23532 6196
rect 23860 5710 23888 6258
rect 23940 5772 23992 5778
rect 23940 5714 23992 5720
rect 23664 5704 23716 5710
rect 23664 5646 23716 5652
rect 23756 5704 23808 5710
rect 23756 5646 23808 5652
rect 23848 5704 23900 5710
rect 23848 5646 23900 5652
rect 22928 5364 22980 5370
rect 22928 5306 22980 5312
rect 23204 5364 23256 5370
rect 23204 5306 23256 5312
rect 22940 5234 22968 5306
rect 22928 5228 22980 5234
rect 22928 5170 22980 5176
rect 23020 5092 23072 5098
rect 23020 5034 23072 5040
rect 22744 4616 22796 4622
rect 22744 4558 22796 4564
rect 22652 4480 22704 4486
rect 22652 4422 22704 4428
rect 22664 4146 22692 4422
rect 22652 4140 22704 4146
rect 22652 4082 22704 4088
rect 22756 3738 22784 4558
rect 22836 4548 22888 4554
rect 22836 4490 22888 4496
rect 22848 4146 22876 4490
rect 22928 4480 22980 4486
rect 22928 4422 22980 4428
rect 22836 4140 22888 4146
rect 22836 4082 22888 4088
rect 22940 4010 22968 4422
rect 23032 4282 23060 5034
rect 23296 4820 23348 4826
rect 23296 4762 23348 4768
rect 23308 4570 23336 4762
rect 23112 4548 23164 4554
rect 23112 4490 23164 4496
rect 23216 4542 23336 4570
rect 23020 4276 23072 4282
rect 23020 4218 23072 4224
rect 23124 4146 23152 4490
rect 23020 4140 23072 4146
rect 23020 4082 23072 4088
rect 23112 4140 23164 4146
rect 23112 4082 23164 4088
rect 22928 4004 22980 4010
rect 22928 3946 22980 3952
rect 23032 3738 23060 4082
rect 22744 3732 22796 3738
rect 22744 3674 22796 3680
rect 23020 3732 23072 3738
rect 23020 3674 23072 3680
rect 23124 3466 23152 4082
rect 22560 3460 22612 3466
rect 22560 3402 22612 3408
rect 23112 3460 23164 3466
rect 23112 3402 23164 3408
rect 21824 3392 21876 3398
rect 21824 3334 21876 3340
rect 22652 3392 22704 3398
rect 22652 3334 22704 3340
rect 21732 3120 21784 3126
rect 21732 3062 21784 3068
rect 21836 3058 21864 3334
rect 21824 3052 21876 3058
rect 21824 2994 21876 3000
rect 22100 2984 22152 2990
rect 22100 2926 22152 2932
rect 21456 2916 21508 2922
rect 21456 2858 21508 2864
rect 22112 2650 22140 2926
rect 21180 2644 21232 2650
rect 21180 2586 21232 2592
rect 21272 2644 21324 2650
rect 21272 2586 21324 2592
rect 22100 2644 22152 2650
rect 22100 2586 22152 2592
rect 22664 2514 22692 3334
rect 22652 2508 22704 2514
rect 22652 2450 22704 2456
rect 23124 2446 23152 3402
rect 23216 2802 23244 4542
rect 23296 4480 23348 4486
rect 23296 4422 23348 4428
rect 23480 4480 23532 4486
rect 23480 4422 23532 4428
rect 23308 3534 23336 4422
rect 23388 3936 23440 3942
rect 23388 3878 23440 3884
rect 23400 3738 23428 3878
rect 23388 3732 23440 3738
rect 23388 3674 23440 3680
rect 23296 3528 23348 3534
rect 23296 3470 23348 3476
rect 23296 3392 23348 3398
rect 23296 3334 23348 3340
rect 23308 2938 23336 3334
rect 23400 3074 23428 3674
rect 23492 3534 23520 4422
rect 23572 4276 23624 4282
rect 23572 4218 23624 4224
rect 23584 4146 23612 4218
rect 23572 4140 23624 4146
rect 23572 4082 23624 4088
rect 23676 3942 23704 5646
rect 23768 5370 23796 5646
rect 23756 5364 23808 5370
rect 23756 5306 23808 5312
rect 23756 5228 23808 5234
rect 23860 5216 23888 5646
rect 23952 5234 23980 5714
rect 23808 5188 23888 5216
rect 23940 5228 23992 5234
rect 23756 5170 23808 5176
rect 23940 5170 23992 5176
rect 23768 5030 23796 5170
rect 23756 5024 23808 5030
rect 23756 4966 23808 4972
rect 24044 4826 24072 6258
rect 24216 6248 24268 6254
rect 24216 6190 24268 6196
rect 24492 6248 24544 6254
rect 24492 6190 24544 6196
rect 24584 6248 24636 6254
rect 24584 6190 24636 6196
rect 24032 4820 24084 4826
rect 24032 4762 24084 4768
rect 24044 4282 24072 4762
rect 24228 4690 24256 6190
rect 24504 5914 24532 6190
rect 24596 5914 24624 6190
rect 24492 5908 24544 5914
rect 24492 5850 24544 5856
rect 24584 5908 24636 5914
rect 24584 5850 24636 5856
rect 24780 5778 24808 6326
rect 24964 5794 24992 6326
rect 25044 6112 25096 6118
rect 25044 6054 25096 6060
rect 25056 5914 25084 6054
rect 25148 5914 25176 6598
rect 25516 6254 25544 6598
rect 25504 6248 25556 6254
rect 25504 6190 25556 6196
rect 25261 6012 25569 6021
rect 25261 6010 25267 6012
rect 25323 6010 25347 6012
rect 25403 6010 25427 6012
rect 25483 6010 25507 6012
rect 25563 6010 25569 6012
rect 25323 5958 25325 6010
rect 25505 5958 25507 6010
rect 25261 5956 25267 5958
rect 25323 5956 25347 5958
rect 25403 5956 25427 5958
rect 25483 5956 25507 5958
rect 25563 5956 25569 5958
rect 25261 5947 25569 5956
rect 25044 5908 25096 5914
rect 25044 5850 25096 5856
rect 25136 5908 25188 5914
rect 25136 5850 25188 5856
rect 24768 5772 24820 5778
rect 24964 5766 25176 5794
rect 24768 5714 24820 5720
rect 24308 5636 24360 5642
rect 24308 5578 24360 5584
rect 24320 5234 24348 5578
rect 24308 5228 24360 5234
rect 24308 5170 24360 5176
rect 24860 5228 24912 5234
rect 24860 5170 24912 5176
rect 24676 5024 24728 5030
rect 24676 4966 24728 4972
rect 24688 4690 24716 4966
rect 24216 4684 24268 4690
rect 24216 4626 24268 4632
rect 24676 4684 24728 4690
rect 24676 4626 24728 4632
rect 24032 4276 24084 4282
rect 24032 4218 24084 4224
rect 23664 3936 23716 3942
rect 23664 3878 23716 3884
rect 23756 3936 23808 3942
rect 23756 3878 23808 3884
rect 23768 3534 23796 3878
rect 24228 3602 24256 4626
rect 24872 4162 24900 5170
rect 25148 4554 25176 5766
rect 25608 5710 25636 6938
rect 25688 6792 25740 6798
rect 25688 6734 25740 6740
rect 25700 5846 25728 6734
rect 25921 6556 26229 6565
rect 25921 6554 25927 6556
rect 25983 6554 26007 6556
rect 26063 6554 26087 6556
rect 26143 6554 26167 6556
rect 26223 6554 26229 6556
rect 25983 6502 25985 6554
rect 26165 6502 26167 6554
rect 25921 6500 25927 6502
rect 25983 6500 26007 6502
rect 26063 6500 26087 6502
rect 26143 6500 26167 6502
rect 26223 6500 26229 6502
rect 25921 6491 26229 6500
rect 28276 6322 28304 7754
rect 28264 6316 28316 6322
rect 28264 6258 28316 6264
rect 28540 6248 28592 6254
rect 28538 6216 28540 6225
rect 28592 6216 28594 6225
rect 28538 6151 28594 6160
rect 25688 5840 25740 5846
rect 25688 5782 25740 5788
rect 25596 5704 25648 5710
rect 25596 5646 25648 5652
rect 25608 5234 25636 5646
rect 25700 5234 25728 5782
rect 25921 5468 26229 5477
rect 25921 5466 25927 5468
rect 25983 5466 26007 5468
rect 26063 5466 26087 5468
rect 26143 5466 26167 5468
rect 26223 5466 26229 5468
rect 25983 5414 25985 5466
rect 26165 5414 26167 5466
rect 25921 5412 25927 5414
rect 25983 5412 26007 5414
rect 26063 5412 26087 5414
rect 26143 5412 26167 5414
rect 26223 5412 26229 5414
rect 25921 5403 26229 5412
rect 25596 5228 25648 5234
rect 25596 5170 25648 5176
rect 25688 5228 25740 5234
rect 25688 5170 25740 5176
rect 26148 5024 26200 5030
rect 26148 4966 26200 4972
rect 25261 4924 25569 4933
rect 25261 4922 25267 4924
rect 25323 4922 25347 4924
rect 25403 4922 25427 4924
rect 25483 4922 25507 4924
rect 25563 4922 25569 4924
rect 25323 4870 25325 4922
rect 25505 4870 25507 4922
rect 25261 4868 25267 4870
rect 25323 4868 25347 4870
rect 25403 4868 25427 4870
rect 25483 4868 25507 4870
rect 25563 4868 25569 4870
rect 25261 4859 25569 4868
rect 26160 4826 26188 4966
rect 26148 4820 26200 4826
rect 26148 4762 26200 4768
rect 24952 4548 25004 4554
rect 24952 4490 25004 4496
rect 25136 4548 25188 4554
rect 25136 4490 25188 4496
rect 24964 4282 24992 4490
rect 24952 4276 25004 4282
rect 24952 4218 25004 4224
rect 24780 4134 24900 4162
rect 24780 4078 24808 4134
rect 24768 4072 24820 4078
rect 24768 4014 24820 4020
rect 24216 3596 24268 3602
rect 24216 3538 24268 3544
rect 23480 3528 23532 3534
rect 23480 3470 23532 3476
rect 23756 3528 23808 3534
rect 23756 3470 23808 3476
rect 25148 3466 25176 4490
rect 25921 4380 26229 4389
rect 25921 4378 25927 4380
rect 25983 4378 26007 4380
rect 26063 4378 26087 4380
rect 26143 4378 26167 4380
rect 26223 4378 26229 4380
rect 25983 4326 25985 4378
rect 26165 4326 26167 4378
rect 25921 4324 25927 4326
rect 25983 4324 26007 4326
rect 26063 4324 26087 4326
rect 26143 4324 26167 4326
rect 26223 4324 26229 4326
rect 25921 4315 26229 4324
rect 26148 4072 26200 4078
rect 26148 4014 26200 4020
rect 25261 3836 25569 3845
rect 25261 3834 25267 3836
rect 25323 3834 25347 3836
rect 25403 3834 25427 3836
rect 25483 3834 25507 3836
rect 25563 3834 25569 3836
rect 25323 3782 25325 3834
rect 25505 3782 25507 3834
rect 25261 3780 25267 3782
rect 25323 3780 25347 3782
rect 25403 3780 25427 3782
rect 25483 3780 25507 3782
rect 25563 3780 25569 3782
rect 25261 3771 25569 3780
rect 26160 3738 26188 4014
rect 26148 3732 26200 3738
rect 26148 3674 26200 3680
rect 25136 3460 25188 3466
rect 25136 3402 25188 3408
rect 23400 3046 23520 3074
rect 25148 3058 25176 3402
rect 25921 3292 26229 3301
rect 25921 3290 25927 3292
rect 25983 3290 26007 3292
rect 26063 3290 26087 3292
rect 26143 3290 26167 3292
rect 26223 3290 26229 3292
rect 25983 3238 25985 3290
rect 26165 3238 26167 3290
rect 25921 3236 25927 3238
rect 25983 3236 26007 3238
rect 26063 3236 26087 3238
rect 26143 3236 26167 3238
rect 26223 3236 26229 3238
rect 25921 3227 26229 3236
rect 23492 2990 23520 3046
rect 25136 3052 25188 3058
rect 25136 2994 25188 3000
rect 23480 2984 23532 2990
rect 23308 2910 23428 2938
rect 23480 2926 23532 2932
rect 23216 2774 23336 2802
rect 23308 2650 23336 2774
rect 23296 2644 23348 2650
rect 23296 2586 23348 2592
rect 23400 2446 23428 2910
rect 23664 2848 23716 2854
rect 23664 2790 23716 2796
rect 23676 2514 23704 2790
rect 25261 2748 25569 2757
rect 25261 2746 25267 2748
rect 25323 2746 25347 2748
rect 25403 2746 25427 2748
rect 25483 2746 25507 2748
rect 25563 2746 25569 2748
rect 25323 2694 25325 2746
rect 25505 2694 25507 2746
rect 25261 2692 25267 2694
rect 25323 2692 25347 2694
rect 25403 2692 25427 2694
rect 25483 2692 25507 2694
rect 25563 2692 25569 2694
rect 25261 2683 25569 2692
rect 23664 2508 23716 2514
rect 23664 2450 23716 2456
rect 19616 2440 19668 2446
rect 19616 2382 19668 2388
rect 20720 2440 20772 2446
rect 20720 2382 20772 2388
rect 20904 2440 20956 2446
rect 20904 2382 20956 2388
rect 23112 2440 23164 2446
rect 23112 2382 23164 2388
rect 23388 2440 23440 2446
rect 23388 2382 23440 2388
rect 27068 2440 27120 2446
rect 27068 2382 27120 2388
rect 18788 2304 18840 2310
rect 18788 2246 18840 2252
rect 18975 2204 19283 2213
rect 18975 2202 18981 2204
rect 19037 2202 19061 2204
rect 19117 2202 19141 2204
rect 19197 2202 19221 2204
rect 19277 2202 19283 2204
rect 19037 2150 19039 2202
rect 19219 2150 19221 2202
rect 18975 2148 18981 2150
rect 19037 2148 19061 2150
rect 19117 2148 19141 2150
rect 19197 2148 19221 2150
rect 19277 2148 19283 2150
rect 18975 2139 19283 2148
rect 25921 2204 26229 2213
rect 25921 2202 25927 2204
rect 25983 2202 26007 2204
rect 26063 2202 26087 2204
rect 26143 2202 26167 2204
rect 26223 2202 26229 2204
rect 25983 2150 25985 2202
rect 26165 2150 26167 2202
rect 25921 2148 25927 2150
rect 25983 2148 26007 2150
rect 26063 2148 26087 2150
rect 26143 2148 26167 2150
rect 26223 2148 26229 2150
rect 25921 2139 26229 2148
rect 27080 800 27108 2382
rect 18 0 74 800
rect 9034 0 9090 800
rect 18050 0 18106 800
rect 27066 0 27122 800
<< via2 >>
rect 4429 27770 4485 27772
rect 4509 27770 4565 27772
rect 4589 27770 4645 27772
rect 4669 27770 4725 27772
rect 4429 27718 4475 27770
rect 4475 27718 4485 27770
rect 4509 27718 4539 27770
rect 4539 27718 4551 27770
rect 4551 27718 4565 27770
rect 4589 27718 4603 27770
rect 4603 27718 4615 27770
rect 4615 27718 4645 27770
rect 4669 27718 4679 27770
rect 4679 27718 4725 27770
rect 4429 27716 4485 27718
rect 4509 27716 4565 27718
rect 4589 27716 4645 27718
rect 4669 27716 4725 27718
rect 1490 27648 1546 27704
rect 11375 27770 11431 27772
rect 11455 27770 11511 27772
rect 11535 27770 11591 27772
rect 11615 27770 11671 27772
rect 11375 27718 11421 27770
rect 11421 27718 11431 27770
rect 11455 27718 11485 27770
rect 11485 27718 11497 27770
rect 11497 27718 11511 27770
rect 11535 27718 11549 27770
rect 11549 27718 11561 27770
rect 11561 27718 11591 27770
rect 11615 27718 11625 27770
rect 11625 27718 11671 27770
rect 11375 27716 11431 27718
rect 11455 27716 11511 27718
rect 11535 27716 11591 27718
rect 11615 27716 11671 27718
rect 18321 27770 18377 27772
rect 18401 27770 18457 27772
rect 18481 27770 18537 27772
rect 18561 27770 18617 27772
rect 18321 27718 18367 27770
rect 18367 27718 18377 27770
rect 18401 27718 18431 27770
rect 18431 27718 18443 27770
rect 18443 27718 18457 27770
rect 18481 27718 18495 27770
rect 18495 27718 18507 27770
rect 18507 27718 18537 27770
rect 18561 27718 18571 27770
rect 18571 27718 18617 27770
rect 18321 27716 18377 27718
rect 18401 27716 18457 27718
rect 18481 27716 18537 27718
rect 18561 27716 18617 27718
rect 5089 27226 5145 27228
rect 5169 27226 5225 27228
rect 5249 27226 5305 27228
rect 5329 27226 5385 27228
rect 5089 27174 5135 27226
rect 5135 27174 5145 27226
rect 5169 27174 5199 27226
rect 5199 27174 5211 27226
rect 5211 27174 5225 27226
rect 5249 27174 5263 27226
rect 5263 27174 5275 27226
rect 5275 27174 5305 27226
rect 5329 27174 5339 27226
rect 5339 27174 5385 27226
rect 5089 27172 5145 27174
rect 5169 27172 5225 27174
rect 5249 27172 5305 27174
rect 5329 27172 5385 27174
rect 12035 27226 12091 27228
rect 12115 27226 12171 27228
rect 12195 27226 12251 27228
rect 12275 27226 12331 27228
rect 12035 27174 12081 27226
rect 12081 27174 12091 27226
rect 12115 27174 12145 27226
rect 12145 27174 12157 27226
rect 12157 27174 12171 27226
rect 12195 27174 12209 27226
rect 12209 27174 12221 27226
rect 12221 27174 12251 27226
rect 12275 27174 12285 27226
rect 12285 27174 12331 27226
rect 12035 27172 12091 27174
rect 12115 27172 12171 27174
rect 12195 27172 12251 27174
rect 12275 27172 12331 27174
rect 4429 26682 4485 26684
rect 4509 26682 4565 26684
rect 4589 26682 4645 26684
rect 4669 26682 4725 26684
rect 4429 26630 4475 26682
rect 4475 26630 4485 26682
rect 4509 26630 4539 26682
rect 4539 26630 4551 26682
rect 4551 26630 4565 26682
rect 4589 26630 4603 26682
rect 4603 26630 4615 26682
rect 4615 26630 4645 26682
rect 4669 26630 4679 26682
rect 4679 26630 4725 26682
rect 4429 26628 4485 26630
rect 4509 26628 4565 26630
rect 4589 26628 4645 26630
rect 4669 26628 4725 26630
rect 11375 26682 11431 26684
rect 11455 26682 11511 26684
rect 11535 26682 11591 26684
rect 11615 26682 11671 26684
rect 11375 26630 11421 26682
rect 11421 26630 11431 26682
rect 11455 26630 11485 26682
rect 11485 26630 11497 26682
rect 11497 26630 11511 26682
rect 11535 26630 11549 26682
rect 11549 26630 11561 26682
rect 11561 26630 11591 26682
rect 11615 26630 11625 26682
rect 11625 26630 11671 26682
rect 11375 26628 11431 26630
rect 11455 26628 11511 26630
rect 11535 26628 11591 26630
rect 11615 26628 11671 26630
rect 5089 26138 5145 26140
rect 5169 26138 5225 26140
rect 5249 26138 5305 26140
rect 5329 26138 5385 26140
rect 5089 26086 5135 26138
rect 5135 26086 5145 26138
rect 5169 26086 5199 26138
rect 5199 26086 5211 26138
rect 5211 26086 5225 26138
rect 5249 26086 5263 26138
rect 5263 26086 5275 26138
rect 5275 26086 5305 26138
rect 5329 26086 5339 26138
rect 5339 26086 5385 26138
rect 5089 26084 5145 26086
rect 5169 26084 5225 26086
rect 5249 26084 5305 26086
rect 5329 26084 5385 26086
rect 12035 26138 12091 26140
rect 12115 26138 12171 26140
rect 12195 26138 12251 26140
rect 12275 26138 12331 26140
rect 12035 26086 12081 26138
rect 12081 26086 12091 26138
rect 12115 26086 12145 26138
rect 12145 26086 12157 26138
rect 12157 26086 12171 26138
rect 12195 26086 12209 26138
rect 12209 26086 12221 26138
rect 12221 26086 12251 26138
rect 12275 26086 12285 26138
rect 12285 26086 12331 26138
rect 12035 26084 12091 26086
rect 12115 26084 12171 26086
rect 12195 26084 12251 26086
rect 12275 26084 12331 26086
rect 4429 25594 4485 25596
rect 4509 25594 4565 25596
rect 4589 25594 4645 25596
rect 4669 25594 4725 25596
rect 4429 25542 4475 25594
rect 4475 25542 4485 25594
rect 4509 25542 4539 25594
rect 4539 25542 4551 25594
rect 4551 25542 4565 25594
rect 4589 25542 4603 25594
rect 4603 25542 4615 25594
rect 4615 25542 4645 25594
rect 4669 25542 4679 25594
rect 4679 25542 4725 25594
rect 4429 25540 4485 25542
rect 4509 25540 4565 25542
rect 4589 25540 4645 25542
rect 4669 25540 4725 25542
rect 11375 25594 11431 25596
rect 11455 25594 11511 25596
rect 11535 25594 11591 25596
rect 11615 25594 11671 25596
rect 11375 25542 11421 25594
rect 11421 25542 11431 25594
rect 11455 25542 11485 25594
rect 11485 25542 11497 25594
rect 11497 25542 11511 25594
rect 11535 25542 11549 25594
rect 11549 25542 11561 25594
rect 11561 25542 11591 25594
rect 11615 25542 11625 25594
rect 11625 25542 11671 25594
rect 11375 25540 11431 25542
rect 11455 25540 11511 25542
rect 11535 25540 11591 25542
rect 11615 25540 11671 25542
rect 5089 25050 5145 25052
rect 5169 25050 5225 25052
rect 5249 25050 5305 25052
rect 5329 25050 5385 25052
rect 5089 24998 5135 25050
rect 5135 24998 5145 25050
rect 5169 24998 5199 25050
rect 5199 24998 5211 25050
rect 5211 24998 5225 25050
rect 5249 24998 5263 25050
rect 5263 24998 5275 25050
rect 5275 24998 5305 25050
rect 5329 24998 5339 25050
rect 5339 24998 5385 25050
rect 5089 24996 5145 24998
rect 5169 24996 5225 24998
rect 5249 24996 5305 24998
rect 5329 24996 5385 24998
rect 12035 25050 12091 25052
rect 12115 25050 12171 25052
rect 12195 25050 12251 25052
rect 12275 25050 12331 25052
rect 12035 24998 12081 25050
rect 12081 24998 12091 25050
rect 12115 24998 12145 25050
rect 12145 24998 12157 25050
rect 12157 24998 12171 25050
rect 12195 24998 12209 25050
rect 12209 24998 12221 25050
rect 12221 24998 12251 25050
rect 12275 24998 12285 25050
rect 12285 24998 12331 25050
rect 12035 24996 12091 24998
rect 12115 24996 12171 24998
rect 12195 24996 12251 24998
rect 12275 24996 12331 24998
rect 4429 24506 4485 24508
rect 4509 24506 4565 24508
rect 4589 24506 4645 24508
rect 4669 24506 4725 24508
rect 4429 24454 4475 24506
rect 4475 24454 4485 24506
rect 4509 24454 4539 24506
rect 4539 24454 4551 24506
rect 4551 24454 4565 24506
rect 4589 24454 4603 24506
rect 4603 24454 4615 24506
rect 4615 24454 4645 24506
rect 4669 24454 4679 24506
rect 4679 24454 4725 24506
rect 4429 24452 4485 24454
rect 4509 24452 4565 24454
rect 4589 24452 4645 24454
rect 4669 24452 4725 24454
rect 11375 24506 11431 24508
rect 11455 24506 11511 24508
rect 11535 24506 11591 24508
rect 11615 24506 11671 24508
rect 11375 24454 11421 24506
rect 11421 24454 11431 24506
rect 11455 24454 11485 24506
rect 11485 24454 11497 24506
rect 11497 24454 11511 24506
rect 11535 24454 11549 24506
rect 11549 24454 11561 24506
rect 11561 24454 11591 24506
rect 11615 24454 11625 24506
rect 11625 24454 11671 24506
rect 11375 24452 11431 24454
rect 11455 24452 11511 24454
rect 11535 24452 11591 24454
rect 11615 24452 11671 24454
rect 5089 23962 5145 23964
rect 5169 23962 5225 23964
rect 5249 23962 5305 23964
rect 5329 23962 5385 23964
rect 5089 23910 5135 23962
rect 5135 23910 5145 23962
rect 5169 23910 5199 23962
rect 5199 23910 5211 23962
rect 5211 23910 5225 23962
rect 5249 23910 5263 23962
rect 5263 23910 5275 23962
rect 5275 23910 5305 23962
rect 5329 23910 5339 23962
rect 5339 23910 5385 23962
rect 5089 23908 5145 23910
rect 5169 23908 5225 23910
rect 5249 23908 5305 23910
rect 5329 23908 5385 23910
rect 12035 23962 12091 23964
rect 12115 23962 12171 23964
rect 12195 23962 12251 23964
rect 12275 23962 12331 23964
rect 12035 23910 12081 23962
rect 12081 23910 12091 23962
rect 12115 23910 12145 23962
rect 12145 23910 12157 23962
rect 12157 23910 12171 23962
rect 12195 23910 12209 23962
rect 12209 23910 12221 23962
rect 12221 23910 12251 23962
rect 12275 23910 12285 23962
rect 12285 23910 12331 23962
rect 12035 23908 12091 23910
rect 12115 23908 12171 23910
rect 12195 23908 12251 23910
rect 12275 23908 12331 23910
rect 4429 23418 4485 23420
rect 4509 23418 4565 23420
rect 4589 23418 4645 23420
rect 4669 23418 4725 23420
rect 4429 23366 4475 23418
rect 4475 23366 4485 23418
rect 4509 23366 4539 23418
rect 4539 23366 4551 23418
rect 4551 23366 4565 23418
rect 4589 23366 4603 23418
rect 4603 23366 4615 23418
rect 4615 23366 4645 23418
rect 4669 23366 4679 23418
rect 4679 23366 4725 23418
rect 4429 23364 4485 23366
rect 4509 23364 4565 23366
rect 4589 23364 4645 23366
rect 4669 23364 4725 23366
rect 11375 23418 11431 23420
rect 11455 23418 11511 23420
rect 11535 23418 11591 23420
rect 11615 23418 11671 23420
rect 11375 23366 11421 23418
rect 11421 23366 11431 23418
rect 11455 23366 11485 23418
rect 11485 23366 11497 23418
rect 11497 23366 11511 23418
rect 11535 23366 11549 23418
rect 11549 23366 11561 23418
rect 11561 23366 11591 23418
rect 11615 23366 11625 23418
rect 11625 23366 11671 23418
rect 11375 23364 11431 23366
rect 11455 23364 11511 23366
rect 11535 23364 11591 23366
rect 11615 23364 11671 23366
rect 5089 22874 5145 22876
rect 5169 22874 5225 22876
rect 5249 22874 5305 22876
rect 5329 22874 5385 22876
rect 5089 22822 5135 22874
rect 5135 22822 5145 22874
rect 5169 22822 5199 22874
rect 5199 22822 5211 22874
rect 5211 22822 5225 22874
rect 5249 22822 5263 22874
rect 5263 22822 5275 22874
rect 5275 22822 5305 22874
rect 5329 22822 5339 22874
rect 5339 22822 5385 22874
rect 5089 22820 5145 22822
rect 5169 22820 5225 22822
rect 5249 22820 5305 22822
rect 5329 22820 5385 22822
rect 12035 22874 12091 22876
rect 12115 22874 12171 22876
rect 12195 22874 12251 22876
rect 12275 22874 12331 22876
rect 12035 22822 12081 22874
rect 12081 22822 12091 22874
rect 12115 22822 12145 22874
rect 12145 22822 12157 22874
rect 12157 22822 12171 22874
rect 12195 22822 12209 22874
rect 12209 22822 12221 22874
rect 12221 22822 12251 22874
rect 12275 22822 12285 22874
rect 12285 22822 12331 22874
rect 12035 22820 12091 22822
rect 12115 22820 12171 22822
rect 12195 22820 12251 22822
rect 12275 22820 12331 22822
rect 4429 22330 4485 22332
rect 4509 22330 4565 22332
rect 4589 22330 4645 22332
rect 4669 22330 4725 22332
rect 4429 22278 4475 22330
rect 4475 22278 4485 22330
rect 4509 22278 4539 22330
rect 4539 22278 4551 22330
rect 4551 22278 4565 22330
rect 4589 22278 4603 22330
rect 4603 22278 4615 22330
rect 4615 22278 4645 22330
rect 4669 22278 4679 22330
rect 4679 22278 4725 22330
rect 4429 22276 4485 22278
rect 4509 22276 4565 22278
rect 4589 22276 4645 22278
rect 4669 22276 4725 22278
rect 11375 22330 11431 22332
rect 11455 22330 11511 22332
rect 11535 22330 11591 22332
rect 11615 22330 11671 22332
rect 11375 22278 11421 22330
rect 11421 22278 11431 22330
rect 11455 22278 11485 22330
rect 11485 22278 11497 22330
rect 11497 22278 11511 22330
rect 11535 22278 11549 22330
rect 11549 22278 11561 22330
rect 11561 22278 11591 22330
rect 11615 22278 11625 22330
rect 11625 22278 11671 22330
rect 11375 22276 11431 22278
rect 11455 22276 11511 22278
rect 11535 22276 11591 22278
rect 11615 22276 11671 22278
rect 5089 21786 5145 21788
rect 5169 21786 5225 21788
rect 5249 21786 5305 21788
rect 5329 21786 5385 21788
rect 5089 21734 5135 21786
rect 5135 21734 5145 21786
rect 5169 21734 5199 21786
rect 5199 21734 5211 21786
rect 5211 21734 5225 21786
rect 5249 21734 5263 21786
rect 5263 21734 5275 21786
rect 5275 21734 5305 21786
rect 5329 21734 5339 21786
rect 5339 21734 5385 21786
rect 5089 21732 5145 21734
rect 5169 21732 5225 21734
rect 5249 21732 5305 21734
rect 5329 21732 5385 21734
rect 12035 21786 12091 21788
rect 12115 21786 12171 21788
rect 12195 21786 12251 21788
rect 12275 21786 12331 21788
rect 12035 21734 12081 21786
rect 12081 21734 12091 21786
rect 12115 21734 12145 21786
rect 12145 21734 12157 21786
rect 12157 21734 12171 21786
rect 12195 21734 12209 21786
rect 12209 21734 12221 21786
rect 12221 21734 12251 21786
rect 12275 21734 12285 21786
rect 12285 21734 12331 21786
rect 12035 21732 12091 21734
rect 12115 21732 12171 21734
rect 12195 21732 12251 21734
rect 12275 21732 12331 21734
rect 4429 21242 4485 21244
rect 4509 21242 4565 21244
rect 4589 21242 4645 21244
rect 4669 21242 4725 21244
rect 4429 21190 4475 21242
rect 4475 21190 4485 21242
rect 4509 21190 4539 21242
rect 4539 21190 4551 21242
rect 4551 21190 4565 21242
rect 4589 21190 4603 21242
rect 4603 21190 4615 21242
rect 4615 21190 4645 21242
rect 4669 21190 4679 21242
rect 4679 21190 4725 21242
rect 4429 21188 4485 21190
rect 4509 21188 4565 21190
rect 4589 21188 4645 21190
rect 4669 21188 4725 21190
rect 11375 21242 11431 21244
rect 11455 21242 11511 21244
rect 11535 21242 11591 21244
rect 11615 21242 11671 21244
rect 11375 21190 11421 21242
rect 11421 21190 11431 21242
rect 11455 21190 11485 21242
rect 11485 21190 11497 21242
rect 11497 21190 11511 21242
rect 11535 21190 11549 21242
rect 11549 21190 11561 21242
rect 11561 21190 11591 21242
rect 11615 21190 11625 21242
rect 11625 21190 11671 21242
rect 11375 21188 11431 21190
rect 11455 21188 11511 21190
rect 11535 21188 11591 21190
rect 11615 21188 11671 21190
rect 5089 20698 5145 20700
rect 5169 20698 5225 20700
rect 5249 20698 5305 20700
rect 5329 20698 5385 20700
rect 5089 20646 5135 20698
rect 5135 20646 5145 20698
rect 5169 20646 5199 20698
rect 5199 20646 5211 20698
rect 5211 20646 5225 20698
rect 5249 20646 5263 20698
rect 5263 20646 5275 20698
rect 5275 20646 5305 20698
rect 5329 20646 5339 20698
rect 5339 20646 5385 20698
rect 5089 20644 5145 20646
rect 5169 20644 5225 20646
rect 5249 20644 5305 20646
rect 5329 20644 5385 20646
rect 12035 20698 12091 20700
rect 12115 20698 12171 20700
rect 12195 20698 12251 20700
rect 12275 20698 12331 20700
rect 12035 20646 12081 20698
rect 12081 20646 12091 20698
rect 12115 20646 12145 20698
rect 12145 20646 12157 20698
rect 12157 20646 12171 20698
rect 12195 20646 12209 20698
rect 12209 20646 12221 20698
rect 12221 20646 12251 20698
rect 12275 20646 12285 20698
rect 12285 20646 12331 20698
rect 12035 20644 12091 20646
rect 12115 20644 12171 20646
rect 12195 20644 12251 20646
rect 12275 20644 12331 20646
rect 4429 20154 4485 20156
rect 4509 20154 4565 20156
rect 4589 20154 4645 20156
rect 4669 20154 4725 20156
rect 4429 20102 4475 20154
rect 4475 20102 4485 20154
rect 4509 20102 4539 20154
rect 4539 20102 4551 20154
rect 4551 20102 4565 20154
rect 4589 20102 4603 20154
rect 4603 20102 4615 20154
rect 4615 20102 4645 20154
rect 4669 20102 4679 20154
rect 4679 20102 4725 20154
rect 4429 20100 4485 20102
rect 4509 20100 4565 20102
rect 4589 20100 4645 20102
rect 4669 20100 4725 20102
rect 11375 20154 11431 20156
rect 11455 20154 11511 20156
rect 11535 20154 11591 20156
rect 11615 20154 11671 20156
rect 11375 20102 11421 20154
rect 11421 20102 11431 20154
rect 11455 20102 11485 20154
rect 11485 20102 11497 20154
rect 11497 20102 11511 20154
rect 11535 20102 11549 20154
rect 11549 20102 11561 20154
rect 11561 20102 11591 20154
rect 11615 20102 11625 20154
rect 11625 20102 11671 20154
rect 11375 20100 11431 20102
rect 11455 20100 11511 20102
rect 11535 20100 11591 20102
rect 11615 20100 11671 20102
rect 5089 19610 5145 19612
rect 5169 19610 5225 19612
rect 5249 19610 5305 19612
rect 5329 19610 5385 19612
rect 5089 19558 5135 19610
rect 5135 19558 5145 19610
rect 5169 19558 5199 19610
rect 5199 19558 5211 19610
rect 5211 19558 5225 19610
rect 5249 19558 5263 19610
rect 5263 19558 5275 19610
rect 5275 19558 5305 19610
rect 5329 19558 5339 19610
rect 5339 19558 5385 19610
rect 5089 19556 5145 19558
rect 5169 19556 5225 19558
rect 5249 19556 5305 19558
rect 5329 19556 5385 19558
rect 12035 19610 12091 19612
rect 12115 19610 12171 19612
rect 12195 19610 12251 19612
rect 12275 19610 12331 19612
rect 12035 19558 12081 19610
rect 12081 19558 12091 19610
rect 12115 19558 12145 19610
rect 12145 19558 12157 19610
rect 12157 19558 12171 19610
rect 12195 19558 12209 19610
rect 12209 19558 12221 19610
rect 12221 19558 12251 19610
rect 12275 19558 12285 19610
rect 12285 19558 12331 19610
rect 12035 19556 12091 19558
rect 12115 19556 12171 19558
rect 12195 19556 12251 19558
rect 12275 19556 12331 19558
rect 4429 19066 4485 19068
rect 4509 19066 4565 19068
rect 4589 19066 4645 19068
rect 4669 19066 4725 19068
rect 4429 19014 4475 19066
rect 4475 19014 4485 19066
rect 4509 19014 4539 19066
rect 4539 19014 4551 19066
rect 4551 19014 4565 19066
rect 4589 19014 4603 19066
rect 4603 19014 4615 19066
rect 4615 19014 4645 19066
rect 4669 19014 4679 19066
rect 4679 19014 4725 19066
rect 4429 19012 4485 19014
rect 4509 19012 4565 19014
rect 4589 19012 4645 19014
rect 4669 19012 4725 19014
rect 11375 19066 11431 19068
rect 11455 19066 11511 19068
rect 11535 19066 11591 19068
rect 11615 19066 11671 19068
rect 11375 19014 11421 19066
rect 11421 19014 11431 19066
rect 11455 19014 11485 19066
rect 11485 19014 11497 19066
rect 11497 19014 11511 19066
rect 11535 19014 11549 19066
rect 11549 19014 11561 19066
rect 11561 19014 11591 19066
rect 11615 19014 11625 19066
rect 11625 19014 11671 19066
rect 11375 19012 11431 19014
rect 11455 19012 11511 19014
rect 11535 19012 11591 19014
rect 11615 19012 11671 19014
rect 5089 18522 5145 18524
rect 5169 18522 5225 18524
rect 5249 18522 5305 18524
rect 5329 18522 5385 18524
rect 5089 18470 5135 18522
rect 5135 18470 5145 18522
rect 5169 18470 5199 18522
rect 5199 18470 5211 18522
rect 5211 18470 5225 18522
rect 5249 18470 5263 18522
rect 5263 18470 5275 18522
rect 5275 18470 5305 18522
rect 5329 18470 5339 18522
rect 5339 18470 5385 18522
rect 5089 18468 5145 18470
rect 5169 18468 5225 18470
rect 5249 18468 5305 18470
rect 5329 18468 5385 18470
rect 12035 18522 12091 18524
rect 12115 18522 12171 18524
rect 12195 18522 12251 18524
rect 12275 18522 12331 18524
rect 12035 18470 12081 18522
rect 12081 18470 12091 18522
rect 12115 18470 12145 18522
rect 12145 18470 12157 18522
rect 12157 18470 12171 18522
rect 12195 18470 12209 18522
rect 12209 18470 12221 18522
rect 12221 18470 12251 18522
rect 12275 18470 12285 18522
rect 12285 18470 12331 18522
rect 12035 18468 12091 18470
rect 12115 18468 12171 18470
rect 12195 18468 12251 18470
rect 12275 18468 12331 18470
rect 938 18400 994 18456
rect 4429 17978 4485 17980
rect 4509 17978 4565 17980
rect 4589 17978 4645 17980
rect 4669 17978 4725 17980
rect 4429 17926 4475 17978
rect 4475 17926 4485 17978
rect 4509 17926 4539 17978
rect 4539 17926 4551 17978
rect 4551 17926 4565 17978
rect 4589 17926 4603 17978
rect 4603 17926 4615 17978
rect 4615 17926 4645 17978
rect 4669 17926 4679 17978
rect 4679 17926 4725 17978
rect 4429 17924 4485 17926
rect 4509 17924 4565 17926
rect 4589 17924 4645 17926
rect 4669 17924 4725 17926
rect 11375 17978 11431 17980
rect 11455 17978 11511 17980
rect 11535 17978 11591 17980
rect 11615 17978 11671 17980
rect 11375 17926 11421 17978
rect 11421 17926 11431 17978
rect 11455 17926 11485 17978
rect 11485 17926 11497 17978
rect 11497 17926 11511 17978
rect 11535 17926 11549 17978
rect 11549 17926 11561 17978
rect 11561 17926 11591 17978
rect 11615 17926 11625 17978
rect 11625 17926 11671 17978
rect 11375 17924 11431 17926
rect 11455 17924 11511 17926
rect 11535 17924 11591 17926
rect 11615 17924 11671 17926
rect 5089 17434 5145 17436
rect 5169 17434 5225 17436
rect 5249 17434 5305 17436
rect 5329 17434 5385 17436
rect 5089 17382 5135 17434
rect 5135 17382 5145 17434
rect 5169 17382 5199 17434
rect 5199 17382 5211 17434
rect 5211 17382 5225 17434
rect 5249 17382 5263 17434
rect 5263 17382 5275 17434
rect 5275 17382 5305 17434
rect 5329 17382 5339 17434
rect 5339 17382 5385 17434
rect 5089 17380 5145 17382
rect 5169 17380 5225 17382
rect 5249 17380 5305 17382
rect 5329 17380 5385 17382
rect 12035 17434 12091 17436
rect 12115 17434 12171 17436
rect 12195 17434 12251 17436
rect 12275 17434 12331 17436
rect 12035 17382 12081 17434
rect 12081 17382 12091 17434
rect 12115 17382 12145 17434
rect 12145 17382 12157 17434
rect 12157 17382 12171 17434
rect 12195 17382 12209 17434
rect 12209 17382 12221 17434
rect 12221 17382 12251 17434
rect 12275 17382 12285 17434
rect 12285 17382 12331 17434
rect 12035 17380 12091 17382
rect 12115 17380 12171 17382
rect 12195 17380 12251 17382
rect 12275 17380 12331 17382
rect 4429 16890 4485 16892
rect 4509 16890 4565 16892
rect 4589 16890 4645 16892
rect 4669 16890 4725 16892
rect 4429 16838 4475 16890
rect 4475 16838 4485 16890
rect 4509 16838 4539 16890
rect 4539 16838 4551 16890
rect 4551 16838 4565 16890
rect 4589 16838 4603 16890
rect 4603 16838 4615 16890
rect 4615 16838 4645 16890
rect 4669 16838 4679 16890
rect 4679 16838 4725 16890
rect 4429 16836 4485 16838
rect 4509 16836 4565 16838
rect 4589 16836 4645 16838
rect 4669 16836 4725 16838
rect 11375 16890 11431 16892
rect 11455 16890 11511 16892
rect 11535 16890 11591 16892
rect 11615 16890 11671 16892
rect 11375 16838 11421 16890
rect 11421 16838 11431 16890
rect 11455 16838 11485 16890
rect 11485 16838 11497 16890
rect 11497 16838 11511 16890
rect 11535 16838 11549 16890
rect 11549 16838 11561 16890
rect 11561 16838 11591 16890
rect 11615 16838 11625 16890
rect 11625 16838 11671 16890
rect 11375 16836 11431 16838
rect 11455 16836 11511 16838
rect 11535 16836 11591 16838
rect 11615 16836 11671 16838
rect 5089 16346 5145 16348
rect 5169 16346 5225 16348
rect 5249 16346 5305 16348
rect 5329 16346 5385 16348
rect 5089 16294 5135 16346
rect 5135 16294 5145 16346
rect 5169 16294 5199 16346
rect 5199 16294 5211 16346
rect 5211 16294 5225 16346
rect 5249 16294 5263 16346
rect 5263 16294 5275 16346
rect 5275 16294 5305 16346
rect 5329 16294 5339 16346
rect 5339 16294 5385 16346
rect 5089 16292 5145 16294
rect 5169 16292 5225 16294
rect 5249 16292 5305 16294
rect 5329 16292 5385 16294
rect 12035 16346 12091 16348
rect 12115 16346 12171 16348
rect 12195 16346 12251 16348
rect 12275 16346 12331 16348
rect 12035 16294 12081 16346
rect 12081 16294 12091 16346
rect 12115 16294 12145 16346
rect 12145 16294 12157 16346
rect 12157 16294 12171 16346
rect 12195 16294 12209 16346
rect 12209 16294 12221 16346
rect 12221 16294 12251 16346
rect 12275 16294 12285 16346
rect 12285 16294 12331 16346
rect 12035 16292 12091 16294
rect 12115 16292 12171 16294
rect 12195 16292 12251 16294
rect 12275 16292 12331 16294
rect 4429 15802 4485 15804
rect 4509 15802 4565 15804
rect 4589 15802 4645 15804
rect 4669 15802 4725 15804
rect 4429 15750 4475 15802
rect 4475 15750 4485 15802
rect 4509 15750 4539 15802
rect 4539 15750 4551 15802
rect 4551 15750 4565 15802
rect 4589 15750 4603 15802
rect 4603 15750 4615 15802
rect 4615 15750 4645 15802
rect 4669 15750 4679 15802
rect 4679 15750 4725 15802
rect 4429 15748 4485 15750
rect 4509 15748 4565 15750
rect 4589 15748 4645 15750
rect 4669 15748 4725 15750
rect 11375 15802 11431 15804
rect 11455 15802 11511 15804
rect 11535 15802 11591 15804
rect 11615 15802 11671 15804
rect 11375 15750 11421 15802
rect 11421 15750 11431 15802
rect 11455 15750 11485 15802
rect 11485 15750 11497 15802
rect 11497 15750 11511 15802
rect 11535 15750 11549 15802
rect 11549 15750 11561 15802
rect 11561 15750 11591 15802
rect 11615 15750 11625 15802
rect 11625 15750 11671 15802
rect 11375 15748 11431 15750
rect 11455 15748 11511 15750
rect 11535 15748 11591 15750
rect 11615 15748 11671 15750
rect 5089 15258 5145 15260
rect 5169 15258 5225 15260
rect 5249 15258 5305 15260
rect 5329 15258 5385 15260
rect 5089 15206 5135 15258
rect 5135 15206 5145 15258
rect 5169 15206 5199 15258
rect 5199 15206 5211 15258
rect 5211 15206 5225 15258
rect 5249 15206 5263 15258
rect 5263 15206 5275 15258
rect 5275 15206 5305 15258
rect 5329 15206 5339 15258
rect 5339 15206 5385 15258
rect 5089 15204 5145 15206
rect 5169 15204 5225 15206
rect 5249 15204 5305 15206
rect 5329 15204 5385 15206
rect 12035 15258 12091 15260
rect 12115 15258 12171 15260
rect 12195 15258 12251 15260
rect 12275 15258 12331 15260
rect 12035 15206 12081 15258
rect 12081 15206 12091 15258
rect 12115 15206 12145 15258
rect 12145 15206 12157 15258
rect 12157 15206 12171 15258
rect 12195 15206 12209 15258
rect 12209 15206 12221 15258
rect 12221 15206 12251 15258
rect 12275 15206 12285 15258
rect 12285 15206 12331 15258
rect 12035 15204 12091 15206
rect 12115 15204 12171 15206
rect 12195 15204 12251 15206
rect 12275 15204 12331 15206
rect 4429 14714 4485 14716
rect 4509 14714 4565 14716
rect 4589 14714 4645 14716
rect 4669 14714 4725 14716
rect 4429 14662 4475 14714
rect 4475 14662 4485 14714
rect 4509 14662 4539 14714
rect 4539 14662 4551 14714
rect 4551 14662 4565 14714
rect 4589 14662 4603 14714
rect 4603 14662 4615 14714
rect 4615 14662 4645 14714
rect 4669 14662 4679 14714
rect 4679 14662 4725 14714
rect 4429 14660 4485 14662
rect 4509 14660 4565 14662
rect 4589 14660 4645 14662
rect 4669 14660 4725 14662
rect 11375 14714 11431 14716
rect 11455 14714 11511 14716
rect 11535 14714 11591 14716
rect 11615 14714 11671 14716
rect 11375 14662 11421 14714
rect 11421 14662 11431 14714
rect 11455 14662 11485 14714
rect 11485 14662 11497 14714
rect 11497 14662 11511 14714
rect 11535 14662 11549 14714
rect 11549 14662 11561 14714
rect 11561 14662 11591 14714
rect 11615 14662 11625 14714
rect 11625 14662 11671 14714
rect 11375 14660 11431 14662
rect 11455 14660 11511 14662
rect 11535 14660 11591 14662
rect 11615 14660 11671 14662
rect 5089 14170 5145 14172
rect 5169 14170 5225 14172
rect 5249 14170 5305 14172
rect 5329 14170 5385 14172
rect 5089 14118 5135 14170
rect 5135 14118 5145 14170
rect 5169 14118 5199 14170
rect 5199 14118 5211 14170
rect 5211 14118 5225 14170
rect 5249 14118 5263 14170
rect 5263 14118 5275 14170
rect 5275 14118 5305 14170
rect 5329 14118 5339 14170
rect 5339 14118 5385 14170
rect 5089 14116 5145 14118
rect 5169 14116 5225 14118
rect 5249 14116 5305 14118
rect 5329 14116 5385 14118
rect 12035 14170 12091 14172
rect 12115 14170 12171 14172
rect 12195 14170 12251 14172
rect 12275 14170 12331 14172
rect 12035 14118 12081 14170
rect 12081 14118 12091 14170
rect 12115 14118 12145 14170
rect 12145 14118 12157 14170
rect 12157 14118 12171 14170
rect 12195 14118 12209 14170
rect 12209 14118 12221 14170
rect 12221 14118 12251 14170
rect 12275 14118 12285 14170
rect 12285 14118 12331 14170
rect 12035 14116 12091 14118
rect 12115 14116 12171 14118
rect 12195 14116 12251 14118
rect 12275 14116 12331 14118
rect 4429 13626 4485 13628
rect 4509 13626 4565 13628
rect 4589 13626 4645 13628
rect 4669 13626 4725 13628
rect 4429 13574 4475 13626
rect 4475 13574 4485 13626
rect 4509 13574 4539 13626
rect 4539 13574 4551 13626
rect 4551 13574 4565 13626
rect 4589 13574 4603 13626
rect 4603 13574 4615 13626
rect 4615 13574 4645 13626
rect 4669 13574 4679 13626
rect 4679 13574 4725 13626
rect 4429 13572 4485 13574
rect 4509 13572 4565 13574
rect 4589 13572 4645 13574
rect 4669 13572 4725 13574
rect 11375 13626 11431 13628
rect 11455 13626 11511 13628
rect 11535 13626 11591 13628
rect 11615 13626 11671 13628
rect 11375 13574 11421 13626
rect 11421 13574 11431 13626
rect 11455 13574 11485 13626
rect 11485 13574 11497 13626
rect 11497 13574 11511 13626
rect 11535 13574 11549 13626
rect 11549 13574 11561 13626
rect 11561 13574 11591 13626
rect 11615 13574 11625 13626
rect 11625 13574 11671 13626
rect 11375 13572 11431 13574
rect 11455 13572 11511 13574
rect 11535 13572 11591 13574
rect 11615 13572 11671 13574
rect 5089 13082 5145 13084
rect 5169 13082 5225 13084
rect 5249 13082 5305 13084
rect 5329 13082 5385 13084
rect 5089 13030 5135 13082
rect 5135 13030 5145 13082
rect 5169 13030 5199 13082
rect 5199 13030 5211 13082
rect 5211 13030 5225 13082
rect 5249 13030 5263 13082
rect 5263 13030 5275 13082
rect 5275 13030 5305 13082
rect 5329 13030 5339 13082
rect 5339 13030 5385 13082
rect 5089 13028 5145 13030
rect 5169 13028 5225 13030
rect 5249 13028 5305 13030
rect 5329 13028 5385 13030
rect 12035 13082 12091 13084
rect 12115 13082 12171 13084
rect 12195 13082 12251 13084
rect 12275 13082 12331 13084
rect 12035 13030 12081 13082
rect 12081 13030 12091 13082
rect 12115 13030 12145 13082
rect 12145 13030 12157 13082
rect 12157 13030 12171 13082
rect 12195 13030 12209 13082
rect 12209 13030 12221 13082
rect 12221 13030 12251 13082
rect 12275 13030 12285 13082
rect 12285 13030 12331 13082
rect 12035 13028 12091 13030
rect 12115 13028 12171 13030
rect 12195 13028 12251 13030
rect 12275 13028 12331 13030
rect 4429 12538 4485 12540
rect 4509 12538 4565 12540
rect 4589 12538 4645 12540
rect 4669 12538 4725 12540
rect 4429 12486 4475 12538
rect 4475 12486 4485 12538
rect 4509 12486 4539 12538
rect 4539 12486 4551 12538
rect 4551 12486 4565 12538
rect 4589 12486 4603 12538
rect 4603 12486 4615 12538
rect 4615 12486 4645 12538
rect 4669 12486 4679 12538
rect 4679 12486 4725 12538
rect 4429 12484 4485 12486
rect 4509 12484 4565 12486
rect 4589 12484 4645 12486
rect 4669 12484 4725 12486
rect 11375 12538 11431 12540
rect 11455 12538 11511 12540
rect 11535 12538 11591 12540
rect 11615 12538 11671 12540
rect 11375 12486 11421 12538
rect 11421 12486 11431 12538
rect 11455 12486 11485 12538
rect 11485 12486 11497 12538
rect 11497 12486 11511 12538
rect 11535 12486 11549 12538
rect 11549 12486 11561 12538
rect 11561 12486 11591 12538
rect 11615 12486 11625 12538
rect 11625 12486 11671 12538
rect 11375 12484 11431 12486
rect 11455 12484 11511 12486
rect 11535 12484 11591 12486
rect 11615 12484 11671 12486
rect 5089 11994 5145 11996
rect 5169 11994 5225 11996
rect 5249 11994 5305 11996
rect 5329 11994 5385 11996
rect 5089 11942 5135 11994
rect 5135 11942 5145 11994
rect 5169 11942 5199 11994
rect 5199 11942 5211 11994
rect 5211 11942 5225 11994
rect 5249 11942 5263 11994
rect 5263 11942 5275 11994
rect 5275 11942 5305 11994
rect 5329 11942 5339 11994
rect 5339 11942 5385 11994
rect 5089 11940 5145 11942
rect 5169 11940 5225 11942
rect 5249 11940 5305 11942
rect 5329 11940 5385 11942
rect 12035 11994 12091 11996
rect 12115 11994 12171 11996
rect 12195 11994 12251 11996
rect 12275 11994 12331 11996
rect 12035 11942 12081 11994
rect 12081 11942 12091 11994
rect 12115 11942 12145 11994
rect 12145 11942 12157 11994
rect 12157 11942 12171 11994
rect 12195 11942 12209 11994
rect 12209 11942 12221 11994
rect 12221 11942 12251 11994
rect 12275 11942 12285 11994
rect 12285 11942 12331 11994
rect 12035 11940 12091 11942
rect 12115 11940 12171 11942
rect 12195 11940 12251 11942
rect 12275 11940 12331 11942
rect 4429 11450 4485 11452
rect 4509 11450 4565 11452
rect 4589 11450 4645 11452
rect 4669 11450 4725 11452
rect 4429 11398 4475 11450
rect 4475 11398 4485 11450
rect 4509 11398 4539 11450
rect 4539 11398 4551 11450
rect 4551 11398 4565 11450
rect 4589 11398 4603 11450
rect 4603 11398 4615 11450
rect 4615 11398 4645 11450
rect 4669 11398 4679 11450
rect 4679 11398 4725 11450
rect 4429 11396 4485 11398
rect 4509 11396 4565 11398
rect 4589 11396 4645 11398
rect 4669 11396 4725 11398
rect 11375 11450 11431 11452
rect 11455 11450 11511 11452
rect 11535 11450 11591 11452
rect 11615 11450 11671 11452
rect 11375 11398 11421 11450
rect 11421 11398 11431 11450
rect 11455 11398 11485 11450
rect 11485 11398 11497 11450
rect 11497 11398 11511 11450
rect 11535 11398 11549 11450
rect 11549 11398 11561 11450
rect 11561 11398 11591 11450
rect 11615 11398 11625 11450
rect 11625 11398 11671 11450
rect 11375 11396 11431 11398
rect 11455 11396 11511 11398
rect 11535 11396 11591 11398
rect 11615 11396 11671 11398
rect 5089 10906 5145 10908
rect 5169 10906 5225 10908
rect 5249 10906 5305 10908
rect 5329 10906 5385 10908
rect 5089 10854 5135 10906
rect 5135 10854 5145 10906
rect 5169 10854 5199 10906
rect 5199 10854 5211 10906
rect 5211 10854 5225 10906
rect 5249 10854 5263 10906
rect 5263 10854 5275 10906
rect 5275 10854 5305 10906
rect 5329 10854 5339 10906
rect 5339 10854 5385 10906
rect 5089 10852 5145 10854
rect 5169 10852 5225 10854
rect 5249 10852 5305 10854
rect 5329 10852 5385 10854
rect 12035 10906 12091 10908
rect 12115 10906 12171 10908
rect 12195 10906 12251 10908
rect 12275 10906 12331 10908
rect 12035 10854 12081 10906
rect 12081 10854 12091 10906
rect 12115 10854 12145 10906
rect 12145 10854 12157 10906
rect 12157 10854 12171 10906
rect 12195 10854 12209 10906
rect 12209 10854 12221 10906
rect 12221 10854 12251 10906
rect 12275 10854 12285 10906
rect 12285 10854 12331 10906
rect 12035 10852 12091 10854
rect 12115 10852 12171 10854
rect 12195 10852 12251 10854
rect 12275 10852 12331 10854
rect 4429 10362 4485 10364
rect 4509 10362 4565 10364
rect 4589 10362 4645 10364
rect 4669 10362 4725 10364
rect 4429 10310 4475 10362
rect 4475 10310 4485 10362
rect 4509 10310 4539 10362
rect 4539 10310 4551 10362
rect 4551 10310 4565 10362
rect 4589 10310 4603 10362
rect 4603 10310 4615 10362
rect 4615 10310 4645 10362
rect 4669 10310 4679 10362
rect 4679 10310 4725 10362
rect 4429 10308 4485 10310
rect 4509 10308 4565 10310
rect 4589 10308 4645 10310
rect 4669 10308 4725 10310
rect 11375 10362 11431 10364
rect 11455 10362 11511 10364
rect 11535 10362 11591 10364
rect 11615 10362 11671 10364
rect 11375 10310 11421 10362
rect 11421 10310 11431 10362
rect 11455 10310 11485 10362
rect 11485 10310 11497 10362
rect 11497 10310 11511 10362
rect 11535 10310 11549 10362
rect 11549 10310 11561 10362
rect 11561 10310 11591 10362
rect 11615 10310 11625 10362
rect 11625 10310 11671 10362
rect 11375 10308 11431 10310
rect 11455 10308 11511 10310
rect 11535 10308 11591 10310
rect 11615 10308 11671 10310
rect 5089 9818 5145 9820
rect 5169 9818 5225 9820
rect 5249 9818 5305 9820
rect 5329 9818 5385 9820
rect 5089 9766 5135 9818
rect 5135 9766 5145 9818
rect 5169 9766 5199 9818
rect 5199 9766 5211 9818
rect 5211 9766 5225 9818
rect 5249 9766 5263 9818
rect 5263 9766 5275 9818
rect 5275 9766 5305 9818
rect 5329 9766 5339 9818
rect 5339 9766 5385 9818
rect 5089 9764 5145 9766
rect 5169 9764 5225 9766
rect 5249 9764 5305 9766
rect 5329 9764 5385 9766
rect 12035 9818 12091 9820
rect 12115 9818 12171 9820
rect 12195 9818 12251 9820
rect 12275 9818 12331 9820
rect 12035 9766 12081 9818
rect 12081 9766 12091 9818
rect 12115 9766 12145 9818
rect 12145 9766 12157 9818
rect 12157 9766 12171 9818
rect 12195 9766 12209 9818
rect 12209 9766 12221 9818
rect 12221 9766 12251 9818
rect 12275 9766 12285 9818
rect 12285 9766 12331 9818
rect 12035 9764 12091 9766
rect 12115 9764 12171 9766
rect 12195 9764 12251 9766
rect 12275 9764 12331 9766
rect 4429 9274 4485 9276
rect 4509 9274 4565 9276
rect 4589 9274 4645 9276
rect 4669 9274 4725 9276
rect 4429 9222 4475 9274
rect 4475 9222 4485 9274
rect 4509 9222 4539 9274
rect 4539 9222 4551 9274
rect 4551 9222 4565 9274
rect 4589 9222 4603 9274
rect 4603 9222 4615 9274
rect 4615 9222 4645 9274
rect 4669 9222 4679 9274
rect 4679 9222 4725 9274
rect 4429 9220 4485 9222
rect 4509 9220 4565 9222
rect 4589 9220 4645 9222
rect 4669 9220 4725 9222
rect 11375 9274 11431 9276
rect 11455 9274 11511 9276
rect 11535 9274 11591 9276
rect 11615 9274 11671 9276
rect 11375 9222 11421 9274
rect 11421 9222 11431 9274
rect 11455 9222 11485 9274
rect 11485 9222 11497 9274
rect 11497 9222 11511 9274
rect 11535 9222 11549 9274
rect 11549 9222 11561 9274
rect 11561 9222 11591 9274
rect 11615 9222 11625 9274
rect 11625 9222 11671 9274
rect 11375 9220 11431 9222
rect 11455 9220 11511 9222
rect 11535 9220 11591 9222
rect 11615 9220 11671 9222
rect 938 8916 940 8936
rect 940 8916 992 8936
rect 992 8916 994 8936
rect 938 8880 994 8916
rect 5089 8730 5145 8732
rect 5169 8730 5225 8732
rect 5249 8730 5305 8732
rect 5329 8730 5385 8732
rect 5089 8678 5135 8730
rect 5135 8678 5145 8730
rect 5169 8678 5199 8730
rect 5199 8678 5211 8730
rect 5211 8678 5225 8730
rect 5249 8678 5263 8730
rect 5263 8678 5275 8730
rect 5275 8678 5305 8730
rect 5329 8678 5339 8730
rect 5339 8678 5385 8730
rect 5089 8676 5145 8678
rect 5169 8676 5225 8678
rect 5249 8676 5305 8678
rect 5329 8676 5385 8678
rect 12035 8730 12091 8732
rect 12115 8730 12171 8732
rect 12195 8730 12251 8732
rect 12275 8730 12331 8732
rect 12035 8678 12081 8730
rect 12081 8678 12091 8730
rect 12115 8678 12145 8730
rect 12145 8678 12157 8730
rect 12157 8678 12171 8730
rect 12195 8678 12209 8730
rect 12209 8678 12221 8730
rect 12221 8678 12251 8730
rect 12275 8678 12285 8730
rect 12285 8678 12331 8730
rect 12035 8676 12091 8678
rect 12115 8676 12171 8678
rect 12195 8676 12251 8678
rect 12275 8676 12331 8678
rect 4429 8186 4485 8188
rect 4509 8186 4565 8188
rect 4589 8186 4645 8188
rect 4669 8186 4725 8188
rect 4429 8134 4475 8186
rect 4475 8134 4485 8186
rect 4509 8134 4539 8186
rect 4539 8134 4551 8186
rect 4551 8134 4565 8186
rect 4589 8134 4603 8186
rect 4603 8134 4615 8186
rect 4615 8134 4645 8186
rect 4669 8134 4679 8186
rect 4679 8134 4725 8186
rect 4429 8132 4485 8134
rect 4509 8132 4565 8134
rect 4589 8132 4645 8134
rect 4669 8132 4725 8134
rect 11375 8186 11431 8188
rect 11455 8186 11511 8188
rect 11535 8186 11591 8188
rect 11615 8186 11671 8188
rect 11375 8134 11421 8186
rect 11421 8134 11431 8186
rect 11455 8134 11485 8186
rect 11485 8134 11497 8186
rect 11497 8134 11511 8186
rect 11535 8134 11549 8186
rect 11549 8134 11561 8186
rect 11561 8134 11591 8186
rect 11615 8134 11625 8186
rect 11625 8134 11671 8186
rect 11375 8132 11431 8134
rect 11455 8132 11511 8134
rect 11535 8132 11591 8134
rect 11615 8132 11671 8134
rect 5089 7642 5145 7644
rect 5169 7642 5225 7644
rect 5249 7642 5305 7644
rect 5329 7642 5385 7644
rect 5089 7590 5135 7642
rect 5135 7590 5145 7642
rect 5169 7590 5199 7642
rect 5199 7590 5211 7642
rect 5211 7590 5225 7642
rect 5249 7590 5263 7642
rect 5263 7590 5275 7642
rect 5275 7590 5305 7642
rect 5329 7590 5339 7642
rect 5339 7590 5385 7642
rect 5089 7588 5145 7590
rect 5169 7588 5225 7590
rect 5249 7588 5305 7590
rect 5329 7588 5385 7590
rect 12035 7642 12091 7644
rect 12115 7642 12171 7644
rect 12195 7642 12251 7644
rect 12275 7642 12331 7644
rect 12035 7590 12081 7642
rect 12081 7590 12091 7642
rect 12115 7590 12145 7642
rect 12145 7590 12157 7642
rect 12157 7590 12171 7642
rect 12195 7590 12209 7642
rect 12209 7590 12221 7642
rect 12221 7590 12251 7642
rect 12275 7590 12285 7642
rect 12285 7590 12331 7642
rect 12035 7588 12091 7590
rect 12115 7588 12171 7590
rect 12195 7588 12251 7590
rect 12275 7588 12331 7590
rect 4429 7098 4485 7100
rect 4509 7098 4565 7100
rect 4589 7098 4645 7100
rect 4669 7098 4725 7100
rect 4429 7046 4475 7098
rect 4475 7046 4485 7098
rect 4509 7046 4539 7098
rect 4539 7046 4551 7098
rect 4551 7046 4565 7098
rect 4589 7046 4603 7098
rect 4603 7046 4615 7098
rect 4615 7046 4645 7098
rect 4669 7046 4679 7098
rect 4679 7046 4725 7098
rect 4429 7044 4485 7046
rect 4509 7044 4565 7046
rect 4589 7044 4645 7046
rect 4669 7044 4725 7046
rect 11375 7098 11431 7100
rect 11455 7098 11511 7100
rect 11535 7098 11591 7100
rect 11615 7098 11671 7100
rect 11375 7046 11421 7098
rect 11421 7046 11431 7098
rect 11455 7046 11485 7098
rect 11485 7046 11497 7098
rect 11497 7046 11511 7098
rect 11535 7046 11549 7098
rect 11549 7046 11561 7098
rect 11561 7046 11591 7098
rect 11615 7046 11625 7098
rect 11625 7046 11671 7098
rect 11375 7044 11431 7046
rect 11455 7044 11511 7046
rect 11535 7044 11591 7046
rect 11615 7044 11671 7046
rect 5089 6554 5145 6556
rect 5169 6554 5225 6556
rect 5249 6554 5305 6556
rect 5329 6554 5385 6556
rect 5089 6502 5135 6554
rect 5135 6502 5145 6554
rect 5169 6502 5199 6554
rect 5199 6502 5211 6554
rect 5211 6502 5225 6554
rect 5249 6502 5263 6554
rect 5263 6502 5275 6554
rect 5275 6502 5305 6554
rect 5329 6502 5339 6554
rect 5339 6502 5385 6554
rect 5089 6500 5145 6502
rect 5169 6500 5225 6502
rect 5249 6500 5305 6502
rect 5329 6500 5385 6502
rect 12035 6554 12091 6556
rect 12115 6554 12171 6556
rect 12195 6554 12251 6556
rect 12275 6554 12331 6556
rect 12035 6502 12081 6554
rect 12081 6502 12091 6554
rect 12115 6502 12145 6554
rect 12145 6502 12157 6554
rect 12157 6502 12171 6554
rect 12195 6502 12209 6554
rect 12209 6502 12221 6554
rect 12221 6502 12251 6554
rect 12275 6502 12285 6554
rect 12285 6502 12331 6554
rect 12035 6500 12091 6502
rect 12115 6500 12171 6502
rect 12195 6500 12251 6502
rect 12275 6500 12331 6502
rect 4429 6010 4485 6012
rect 4509 6010 4565 6012
rect 4589 6010 4645 6012
rect 4669 6010 4725 6012
rect 4429 5958 4475 6010
rect 4475 5958 4485 6010
rect 4509 5958 4539 6010
rect 4539 5958 4551 6010
rect 4551 5958 4565 6010
rect 4589 5958 4603 6010
rect 4603 5958 4615 6010
rect 4615 5958 4645 6010
rect 4669 5958 4679 6010
rect 4679 5958 4725 6010
rect 4429 5956 4485 5958
rect 4509 5956 4565 5958
rect 4589 5956 4645 5958
rect 4669 5956 4725 5958
rect 11375 6010 11431 6012
rect 11455 6010 11511 6012
rect 11535 6010 11591 6012
rect 11615 6010 11671 6012
rect 11375 5958 11421 6010
rect 11421 5958 11431 6010
rect 11455 5958 11485 6010
rect 11485 5958 11497 6010
rect 11497 5958 11511 6010
rect 11535 5958 11549 6010
rect 11549 5958 11561 6010
rect 11561 5958 11591 6010
rect 11615 5958 11625 6010
rect 11625 5958 11671 6010
rect 11375 5956 11431 5958
rect 11455 5956 11511 5958
rect 11535 5956 11591 5958
rect 11615 5956 11671 5958
rect 5089 5466 5145 5468
rect 5169 5466 5225 5468
rect 5249 5466 5305 5468
rect 5329 5466 5385 5468
rect 5089 5414 5135 5466
rect 5135 5414 5145 5466
rect 5169 5414 5199 5466
rect 5199 5414 5211 5466
rect 5211 5414 5225 5466
rect 5249 5414 5263 5466
rect 5263 5414 5275 5466
rect 5275 5414 5305 5466
rect 5329 5414 5339 5466
rect 5339 5414 5385 5466
rect 5089 5412 5145 5414
rect 5169 5412 5225 5414
rect 5249 5412 5305 5414
rect 5329 5412 5385 5414
rect 12035 5466 12091 5468
rect 12115 5466 12171 5468
rect 12195 5466 12251 5468
rect 12275 5466 12331 5468
rect 12035 5414 12081 5466
rect 12081 5414 12091 5466
rect 12115 5414 12145 5466
rect 12145 5414 12157 5466
rect 12157 5414 12171 5466
rect 12195 5414 12209 5466
rect 12209 5414 12221 5466
rect 12221 5414 12251 5466
rect 12275 5414 12285 5466
rect 12285 5414 12331 5466
rect 12035 5412 12091 5414
rect 12115 5412 12171 5414
rect 12195 5412 12251 5414
rect 12275 5412 12331 5414
rect 4429 4922 4485 4924
rect 4509 4922 4565 4924
rect 4589 4922 4645 4924
rect 4669 4922 4725 4924
rect 4429 4870 4475 4922
rect 4475 4870 4485 4922
rect 4509 4870 4539 4922
rect 4539 4870 4551 4922
rect 4551 4870 4565 4922
rect 4589 4870 4603 4922
rect 4603 4870 4615 4922
rect 4615 4870 4645 4922
rect 4669 4870 4679 4922
rect 4679 4870 4725 4922
rect 4429 4868 4485 4870
rect 4509 4868 4565 4870
rect 4589 4868 4645 4870
rect 4669 4868 4725 4870
rect 11375 4922 11431 4924
rect 11455 4922 11511 4924
rect 11535 4922 11591 4924
rect 11615 4922 11671 4924
rect 11375 4870 11421 4922
rect 11421 4870 11431 4922
rect 11455 4870 11485 4922
rect 11485 4870 11497 4922
rect 11497 4870 11511 4922
rect 11535 4870 11549 4922
rect 11549 4870 11561 4922
rect 11561 4870 11591 4922
rect 11615 4870 11625 4922
rect 11625 4870 11671 4922
rect 11375 4868 11431 4870
rect 11455 4868 11511 4870
rect 11535 4868 11591 4870
rect 11615 4868 11671 4870
rect 5089 4378 5145 4380
rect 5169 4378 5225 4380
rect 5249 4378 5305 4380
rect 5329 4378 5385 4380
rect 5089 4326 5135 4378
rect 5135 4326 5145 4378
rect 5169 4326 5199 4378
rect 5199 4326 5211 4378
rect 5211 4326 5225 4378
rect 5249 4326 5263 4378
rect 5263 4326 5275 4378
rect 5275 4326 5305 4378
rect 5329 4326 5339 4378
rect 5339 4326 5385 4378
rect 5089 4324 5145 4326
rect 5169 4324 5225 4326
rect 5249 4324 5305 4326
rect 5329 4324 5385 4326
rect 12035 4378 12091 4380
rect 12115 4378 12171 4380
rect 12195 4378 12251 4380
rect 12275 4378 12331 4380
rect 12035 4326 12081 4378
rect 12081 4326 12091 4378
rect 12115 4326 12145 4378
rect 12145 4326 12157 4378
rect 12157 4326 12171 4378
rect 12195 4326 12209 4378
rect 12209 4326 12221 4378
rect 12221 4326 12251 4378
rect 12275 4326 12285 4378
rect 12285 4326 12331 4378
rect 12035 4324 12091 4326
rect 12115 4324 12171 4326
rect 12195 4324 12251 4326
rect 12275 4324 12331 4326
rect 4429 3834 4485 3836
rect 4509 3834 4565 3836
rect 4589 3834 4645 3836
rect 4669 3834 4725 3836
rect 4429 3782 4475 3834
rect 4475 3782 4485 3834
rect 4509 3782 4539 3834
rect 4539 3782 4551 3834
rect 4551 3782 4565 3834
rect 4589 3782 4603 3834
rect 4603 3782 4615 3834
rect 4615 3782 4645 3834
rect 4669 3782 4679 3834
rect 4679 3782 4725 3834
rect 4429 3780 4485 3782
rect 4509 3780 4565 3782
rect 4589 3780 4645 3782
rect 4669 3780 4725 3782
rect 11375 3834 11431 3836
rect 11455 3834 11511 3836
rect 11535 3834 11591 3836
rect 11615 3834 11671 3836
rect 11375 3782 11421 3834
rect 11421 3782 11431 3834
rect 11455 3782 11485 3834
rect 11485 3782 11497 3834
rect 11497 3782 11511 3834
rect 11535 3782 11549 3834
rect 11549 3782 11561 3834
rect 11561 3782 11591 3834
rect 11615 3782 11625 3834
rect 11625 3782 11671 3834
rect 11375 3780 11431 3782
rect 11455 3780 11511 3782
rect 11535 3780 11591 3782
rect 11615 3780 11671 3782
rect 5089 3290 5145 3292
rect 5169 3290 5225 3292
rect 5249 3290 5305 3292
rect 5329 3290 5385 3292
rect 5089 3238 5135 3290
rect 5135 3238 5145 3290
rect 5169 3238 5199 3290
rect 5199 3238 5211 3290
rect 5211 3238 5225 3290
rect 5249 3238 5263 3290
rect 5263 3238 5275 3290
rect 5275 3238 5305 3290
rect 5329 3238 5339 3290
rect 5339 3238 5385 3290
rect 5089 3236 5145 3238
rect 5169 3236 5225 3238
rect 5249 3236 5305 3238
rect 5329 3236 5385 3238
rect 12035 3290 12091 3292
rect 12115 3290 12171 3292
rect 12195 3290 12251 3292
rect 12275 3290 12331 3292
rect 12035 3238 12081 3290
rect 12081 3238 12091 3290
rect 12115 3238 12145 3290
rect 12145 3238 12157 3290
rect 12157 3238 12171 3290
rect 12195 3238 12209 3290
rect 12209 3238 12221 3290
rect 12221 3238 12251 3290
rect 12275 3238 12285 3290
rect 12285 3238 12331 3290
rect 12035 3236 12091 3238
rect 12115 3236 12171 3238
rect 12195 3236 12251 3238
rect 12275 3236 12331 3238
rect 4429 2746 4485 2748
rect 4509 2746 4565 2748
rect 4589 2746 4645 2748
rect 4669 2746 4725 2748
rect 4429 2694 4475 2746
rect 4475 2694 4485 2746
rect 4509 2694 4539 2746
rect 4539 2694 4551 2746
rect 4551 2694 4565 2746
rect 4589 2694 4603 2746
rect 4603 2694 4615 2746
rect 4615 2694 4645 2746
rect 4669 2694 4679 2746
rect 4679 2694 4725 2746
rect 4429 2692 4485 2694
rect 4509 2692 4565 2694
rect 4589 2692 4645 2694
rect 4669 2692 4725 2694
rect 11375 2746 11431 2748
rect 11455 2746 11511 2748
rect 11535 2746 11591 2748
rect 11615 2746 11671 2748
rect 11375 2694 11421 2746
rect 11421 2694 11431 2746
rect 11455 2694 11485 2746
rect 11485 2694 11497 2746
rect 11497 2694 11511 2746
rect 11535 2694 11549 2746
rect 11549 2694 11561 2746
rect 11561 2694 11591 2746
rect 11615 2694 11625 2746
rect 11625 2694 11671 2746
rect 11375 2692 11431 2694
rect 11455 2692 11511 2694
rect 11535 2692 11591 2694
rect 11615 2692 11671 2694
rect 18981 27226 19037 27228
rect 19061 27226 19117 27228
rect 19141 27226 19197 27228
rect 19221 27226 19277 27228
rect 18981 27174 19027 27226
rect 19027 27174 19037 27226
rect 19061 27174 19091 27226
rect 19091 27174 19103 27226
rect 19103 27174 19117 27226
rect 19141 27174 19155 27226
rect 19155 27174 19167 27226
rect 19167 27174 19197 27226
rect 19221 27174 19231 27226
rect 19231 27174 19277 27226
rect 18981 27172 19037 27174
rect 19061 27172 19117 27174
rect 19141 27172 19197 27174
rect 19221 27172 19277 27174
rect 18321 26682 18377 26684
rect 18401 26682 18457 26684
rect 18481 26682 18537 26684
rect 18561 26682 18617 26684
rect 18321 26630 18367 26682
rect 18367 26630 18377 26682
rect 18401 26630 18431 26682
rect 18431 26630 18443 26682
rect 18443 26630 18457 26682
rect 18481 26630 18495 26682
rect 18495 26630 18507 26682
rect 18507 26630 18537 26682
rect 18561 26630 18571 26682
rect 18571 26630 18617 26682
rect 18321 26628 18377 26630
rect 18401 26628 18457 26630
rect 18481 26628 18537 26630
rect 18561 26628 18617 26630
rect 18981 26138 19037 26140
rect 19061 26138 19117 26140
rect 19141 26138 19197 26140
rect 19221 26138 19277 26140
rect 18981 26086 19027 26138
rect 19027 26086 19037 26138
rect 19061 26086 19091 26138
rect 19091 26086 19103 26138
rect 19103 26086 19117 26138
rect 19141 26086 19155 26138
rect 19155 26086 19167 26138
rect 19167 26086 19197 26138
rect 19221 26086 19231 26138
rect 19231 26086 19277 26138
rect 18981 26084 19037 26086
rect 19061 26084 19117 26086
rect 19141 26084 19197 26086
rect 19221 26084 19277 26086
rect 18321 25594 18377 25596
rect 18401 25594 18457 25596
rect 18481 25594 18537 25596
rect 18561 25594 18617 25596
rect 18321 25542 18367 25594
rect 18367 25542 18377 25594
rect 18401 25542 18431 25594
rect 18431 25542 18443 25594
rect 18443 25542 18457 25594
rect 18481 25542 18495 25594
rect 18495 25542 18507 25594
rect 18507 25542 18537 25594
rect 18561 25542 18571 25594
rect 18571 25542 18617 25594
rect 18321 25540 18377 25542
rect 18401 25540 18457 25542
rect 18481 25540 18537 25542
rect 18561 25540 18617 25542
rect 18981 25050 19037 25052
rect 19061 25050 19117 25052
rect 19141 25050 19197 25052
rect 19221 25050 19277 25052
rect 18981 24998 19027 25050
rect 19027 24998 19037 25050
rect 19061 24998 19091 25050
rect 19091 24998 19103 25050
rect 19103 24998 19117 25050
rect 19141 24998 19155 25050
rect 19155 24998 19167 25050
rect 19167 24998 19197 25050
rect 19221 24998 19231 25050
rect 19231 24998 19277 25050
rect 18981 24996 19037 24998
rect 19061 24996 19117 24998
rect 19141 24996 19197 24998
rect 19221 24996 19277 24998
rect 18321 24506 18377 24508
rect 18401 24506 18457 24508
rect 18481 24506 18537 24508
rect 18561 24506 18617 24508
rect 18321 24454 18367 24506
rect 18367 24454 18377 24506
rect 18401 24454 18431 24506
rect 18431 24454 18443 24506
rect 18443 24454 18457 24506
rect 18481 24454 18495 24506
rect 18495 24454 18507 24506
rect 18507 24454 18537 24506
rect 18561 24454 18571 24506
rect 18571 24454 18617 24506
rect 18321 24452 18377 24454
rect 18401 24452 18457 24454
rect 18481 24452 18537 24454
rect 18561 24452 18617 24454
rect 18981 23962 19037 23964
rect 19061 23962 19117 23964
rect 19141 23962 19197 23964
rect 19221 23962 19277 23964
rect 18981 23910 19027 23962
rect 19027 23910 19037 23962
rect 19061 23910 19091 23962
rect 19091 23910 19103 23962
rect 19103 23910 19117 23962
rect 19141 23910 19155 23962
rect 19155 23910 19167 23962
rect 19167 23910 19197 23962
rect 19221 23910 19231 23962
rect 19231 23910 19277 23962
rect 18981 23908 19037 23910
rect 19061 23908 19117 23910
rect 19141 23908 19197 23910
rect 19221 23908 19277 23910
rect 18321 23418 18377 23420
rect 18401 23418 18457 23420
rect 18481 23418 18537 23420
rect 18561 23418 18617 23420
rect 18321 23366 18367 23418
rect 18367 23366 18377 23418
rect 18401 23366 18431 23418
rect 18431 23366 18443 23418
rect 18443 23366 18457 23418
rect 18481 23366 18495 23418
rect 18495 23366 18507 23418
rect 18507 23366 18537 23418
rect 18561 23366 18571 23418
rect 18571 23366 18617 23418
rect 18321 23364 18377 23366
rect 18401 23364 18457 23366
rect 18481 23364 18537 23366
rect 18561 23364 18617 23366
rect 18981 22874 19037 22876
rect 19061 22874 19117 22876
rect 19141 22874 19197 22876
rect 19221 22874 19277 22876
rect 18981 22822 19027 22874
rect 19027 22822 19037 22874
rect 19061 22822 19091 22874
rect 19091 22822 19103 22874
rect 19103 22822 19117 22874
rect 19141 22822 19155 22874
rect 19155 22822 19167 22874
rect 19167 22822 19197 22874
rect 19221 22822 19231 22874
rect 19231 22822 19277 22874
rect 18981 22820 19037 22822
rect 19061 22820 19117 22822
rect 19141 22820 19197 22822
rect 19221 22820 19277 22822
rect 18321 22330 18377 22332
rect 18401 22330 18457 22332
rect 18481 22330 18537 22332
rect 18561 22330 18617 22332
rect 18321 22278 18367 22330
rect 18367 22278 18377 22330
rect 18401 22278 18431 22330
rect 18431 22278 18443 22330
rect 18443 22278 18457 22330
rect 18481 22278 18495 22330
rect 18495 22278 18507 22330
rect 18507 22278 18537 22330
rect 18561 22278 18571 22330
rect 18571 22278 18617 22330
rect 18321 22276 18377 22278
rect 18401 22276 18457 22278
rect 18481 22276 18537 22278
rect 18561 22276 18617 22278
rect 18981 21786 19037 21788
rect 19061 21786 19117 21788
rect 19141 21786 19197 21788
rect 19221 21786 19277 21788
rect 18981 21734 19027 21786
rect 19027 21734 19037 21786
rect 19061 21734 19091 21786
rect 19091 21734 19103 21786
rect 19103 21734 19117 21786
rect 19141 21734 19155 21786
rect 19155 21734 19167 21786
rect 19167 21734 19197 21786
rect 19221 21734 19231 21786
rect 19231 21734 19277 21786
rect 18981 21732 19037 21734
rect 19061 21732 19117 21734
rect 19141 21732 19197 21734
rect 19221 21732 19277 21734
rect 18321 21242 18377 21244
rect 18401 21242 18457 21244
rect 18481 21242 18537 21244
rect 18561 21242 18617 21244
rect 18321 21190 18367 21242
rect 18367 21190 18377 21242
rect 18401 21190 18431 21242
rect 18431 21190 18443 21242
rect 18443 21190 18457 21242
rect 18481 21190 18495 21242
rect 18495 21190 18507 21242
rect 18507 21190 18537 21242
rect 18561 21190 18571 21242
rect 18571 21190 18617 21242
rect 18321 21188 18377 21190
rect 18401 21188 18457 21190
rect 18481 21188 18537 21190
rect 18561 21188 18617 21190
rect 18981 20698 19037 20700
rect 19061 20698 19117 20700
rect 19141 20698 19197 20700
rect 19221 20698 19277 20700
rect 18981 20646 19027 20698
rect 19027 20646 19037 20698
rect 19061 20646 19091 20698
rect 19091 20646 19103 20698
rect 19103 20646 19117 20698
rect 19141 20646 19155 20698
rect 19155 20646 19167 20698
rect 19167 20646 19197 20698
rect 19221 20646 19231 20698
rect 19231 20646 19277 20698
rect 18981 20644 19037 20646
rect 19061 20644 19117 20646
rect 19141 20644 19197 20646
rect 19221 20644 19277 20646
rect 18321 20154 18377 20156
rect 18401 20154 18457 20156
rect 18481 20154 18537 20156
rect 18561 20154 18617 20156
rect 18321 20102 18367 20154
rect 18367 20102 18377 20154
rect 18401 20102 18431 20154
rect 18431 20102 18443 20154
rect 18443 20102 18457 20154
rect 18481 20102 18495 20154
rect 18495 20102 18507 20154
rect 18507 20102 18537 20154
rect 18561 20102 18571 20154
rect 18571 20102 18617 20154
rect 18321 20100 18377 20102
rect 18401 20100 18457 20102
rect 18481 20100 18537 20102
rect 18561 20100 18617 20102
rect 18981 19610 19037 19612
rect 19061 19610 19117 19612
rect 19141 19610 19197 19612
rect 19221 19610 19277 19612
rect 18981 19558 19027 19610
rect 19027 19558 19037 19610
rect 19061 19558 19091 19610
rect 19091 19558 19103 19610
rect 19103 19558 19117 19610
rect 19141 19558 19155 19610
rect 19155 19558 19167 19610
rect 19167 19558 19197 19610
rect 19221 19558 19231 19610
rect 19231 19558 19277 19610
rect 18981 19556 19037 19558
rect 19061 19556 19117 19558
rect 19141 19556 19197 19558
rect 19221 19556 19277 19558
rect 18321 19066 18377 19068
rect 18401 19066 18457 19068
rect 18481 19066 18537 19068
rect 18561 19066 18617 19068
rect 18321 19014 18367 19066
rect 18367 19014 18377 19066
rect 18401 19014 18431 19066
rect 18431 19014 18443 19066
rect 18443 19014 18457 19066
rect 18481 19014 18495 19066
rect 18495 19014 18507 19066
rect 18507 19014 18537 19066
rect 18561 19014 18571 19066
rect 18571 19014 18617 19066
rect 18321 19012 18377 19014
rect 18401 19012 18457 19014
rect 18481 19012 18537 19014
rect 18561 19012 18617 19014
rect 18981 18522 19037 18524
rect 19061 18522 19117 18524
rect 19141 18522 19197 18524
rect 19221 18522 19277 18524
rect 18981 18470 19027 18522
rect 19027 18470 19037 18522
rect 19061 18470 19091 18522
rect 19091 18470 19103 18522
rect 19103 18470 19117 18522
rect 19141 18470 19155 18522
rect 19155 18470 19167 18522
rect 19167 18470 19197 18522
rect 19221 18470 19231 18522
rect 19231 18470 19277 18522
rect 18981 18468 19037 18470
rect 19061 18468 19117 18470
rect 19141 18468 19197 18470
rect 19221 18468 19277 18470
rect 18321 17978 18377 17980
rect 18401 17978 18457 17980
rect 18481 17978 18537 17980
rect 18561 17978 18617 17980
rect 18321 17926 18367 17978
rect 18367 17926 18377 17978
rect 18401 17926 18431 17978
rect 18431 17926 18443 17978
rect 18443 17926 18457 17978
rect 18481 17926 18495 17978
rect 18495 17926 18507 17978
rect 18507 17926 18537 17978
rect 18561 17926 18571 17978
rect 18571 17926 18617 17978
rect 18321 17924 18377 17926
rect 18401 17924 18457 17926
rect 18481 17924 18537 17926
rect 18561 17924 18617 17926
rect 18981 17434 19037 17436
rect 19061 17434 19117 17436
rect 19141 17434 19197 17436
rect 19221 17434 19277 17436
rect 18981 17382 19027 17434
rect 19027 17382 19037 17434
rect 19061 17382 19091 17434
rect 19091 17382 19103 17434
rect 19103 17382 19117 17434
rect 19141 17382 19155 17434
rect 19155 17382 19167 17434
rect 19167 17382 19197 17434
rect 19221 17382 19231 17434
rect 19231 17382 19277 17434
rect 18981 17380 19037 17382
rect 19061 17380 19117 17382
rect 19141 17380 19197 17382
rect 19221 17380 19277 17382
rect 18321 16890 18377 16892
rect 18401 16890 18457 16892
rect 18481 16890 18537 16892
rect 18561 16890 18617 16892
rect 18321 16838 18367 16890
rect 18367 16838 18377 16890
rect 18401 16838 18431 16890
rect 18431 16838 18443 16890
rect 18443 16838 18457 16890
rect 18481 16838 18495 16890
rect 18495 16838 18507 16890
rect 18507 16838 18537 16890
rect 18561 16838 18571 16890
rect 18571 16838 18617 16890
rect 18321 16836 18377 16838
rect 18401 16836 18457 16838
rect 18481 16836 18537 16838
rect 18561 16836 18617 16838
rect 18981 16346 19037 16348
rect 19061 16346 19117 16348
rect 19141 16346 19197 16348
rect 19221 16346 19277 16348
rect 18981 16294 19027 16346
rect 19027 16294 19037 16346
rect 19061 16294 19091 16346
rect 19091 16294 19103 16346
rect 19103 16294 19117 16346
rect 19141 16294 19155 16346
rect 19155 16294 19167 16346
rect 19167 16294 19197 16346
rect 19221 16294 19231 16346
rect 19231 16294 19277 16346
rect 18981 16292 19037 16294
rect 19061 16292 19117 16294
rect 19141 16292 19197 16294
rect 19221 16292 19277 16294
rect 18321 15802 18377 15804
rect 18401 15802 18457 15804
rect 18481 15802 18537 15804
rect 18561 15802 18617 15804
rect 18321 15750 18367 15802
rect 18367 15750 18377 15802
rect 18401 15750 18431 15802
rect 18431 15750 18443 15802
rect 18443 15750 18457 15802
rect 18481 15750 18495 15802
rect 18495 15750 18507 15802
rect 18507 15750 18537 15802
rect 18561 15750 18571 15802
rect 18571 15750 18617 15802
rect 18321 15748 18377 15750
rect 18401 15748 18457 15750
rect 18481 15748 18537 15750
rect 18561 15748 18617 15750
rect 18981 15258 19037 15260
rect 19061 15258 19117 15260
rect 19141 15258 19197 15260
rect 19221 15258 19277 15260
rect 18981 15206 19027 15258
rect 19027 15206 19037 15258
rect 19061 15206 19091 15258
rect 19091 15206 19103 15258
rect 19103 15206 19117 15258
rect 19141 15206 19155 15258
rect 19155 15206 19167 15258
rect 19167 15206 19197 15258
rect 19221 15206 19231 15258
rect 19231 15206 19277 15258
rect 18981 15204 19037 15206
rect 19061 15204 19117 15206
rect 19141 15204 19197 15206
rect 19221 15204 19277 15206
rect 18321 14714 18377 14716
rect 18401 14714 18457 14716
rect 18481 14714 18537 14716
rect 18561 14714 18617 14716
rect 18321 14662 18367 14714
rect 18367 14662 18377 14714
rect 18401 14662 18431 14714
rect 18431 14662 18443 14714
rect 18443 14662 18457 14714
rect 18481 14662 18495 14714
rect 18495 14662 18507 14714
rect 18507 14662 18537 14714
rect 18561 14662 18571 14714
rect 18571 14662 18617 14714
rect 18321 14660 18377 14662
rect 18401 14660 18457 14662
rect 18481 14660 18537 14662
rect 18561 14660 18617 14662
rect 18981 14170 19037 14172
rect 19061 14170 19117 14172
rect 19141 14170 19197 14172
rect 19221 14170 19277 14172
rect 18981 14118 19027 14170
rect 19027 14118 19037 14170
rect 19061 14118 19091 14170
rect 19091 14118 19103 14170
rect 19103 14118 19117 14170
rect 19141 14118 19155 14170
rect 19155 14118 19167 14170
rect 19167 14118 19197 14170
rect 19221 14118 19231 14170
rect 19231 14118 19277 14170
rect 18981 14116 19037 14118
rect 19061 14116 19117 14118
rect 19141 14116 19197 14118
rect 19221 14116 19277 14118
rect 18321 13626 18377 13628
rect 18401 13626 18457 13628
rect 18481 13626 18537 13628
rect 18561 13626 18617 13628
rect 18321 13574 18367 13626
rect 18367 13574 18377 13626
rect 18401 13574 18431 13626
rect 18431 13574 18443 13626
rect 18443 13574 18457 13626
rect 18481 13574 18495 13626
rect 18495 13574 18507 13626
rect 18507 13574 18537 13626
rect 18561 13574 18571 13626
rect 18571 13574 18617 13626
rect 18321 13572 18377 13574
rect 18401 13572 18457 13574
rect 18481 13572 18537 13574
rect 18561 13572 18617 13574
rect 18981 13082 19037 13084
rect 19061 13082 19117 13084
rect 19141 13082 19197 13084
rect 19221 13082 19277 13084
rect 18981 13030 19027 13082
rect 19027 13030 19037 13082
rect 19061 13030 19091 13082
rect 19091 13030 19103 13082
rect 19103 13030 19117 13082
rect 19141 13030 19155 13082
rect 19155 13030 19167 13082
rect 19167 13030 19197 13082
rect 19221 13030 19231 13082
rect 19231 13030 19277 13082
rect 18981 13028 19037 13030
rect 19061 13028 19117 13030
rect 19141 13028 19197 13030
rect 19221 13028 19277 13030
rect 18321 12538 18377 12540
rect 18401 12538 18457 12540
rect 18481 12538 18537 12540
rect 18561 12538 18617 12540
rect 18321 12486 18367 12538
rect 18367 12486 18377 12538
rect 18401 12486 18431 12538
rect 18431 12486 18443 12538
rect 18443 12486 18457 12538
rect 18481 12486 18495 12538
rect 18495 12486 18507 12538
rect 18507 12486 18537 12538
rect 18561 12486 18571 12538
rect 18571 12486 18617 12538
rect 18321 12484 18377 12486
rect 18401 12484 18457 12486
rect 18481 12484 18537 12486
rect 18561 12484 18617 12486
rect 16762 9016 16818 9072
rect 18981 11994 19037 11996
rect 19061 11994 19117 11996
rect 19141 11994 19197 11996
rect 19221 11994 19277 11996
rect 18981 11942 19027 11994
rect 19027 11942 19037 11994
rect 19061 11942 19091 11994
rect 19091 11942 19103 11994
rect 19103 11942 19117 11994
rect 19141 11942 19155 11994
rect 19155 11942 19167 11994
rect 19167 11942 19197 11994
rect 19221 11942 19231 11994
rect 19231 11942 19277 11994
rect 18981 11940 19037 11942
rect 19061 11940 19117 11942
rect 19141 11940 19197 11942
rect 19221 11940 19277 11942
rect 18321 11450 18377 11452
rect 18401 11450 18457 11452
rect 18481 11450 18537 11452
rect 18561 11450 18617 11452
rect 18321 11398 18367 11450
rect 18367 11398 18377 11450
rect 18401 11398 18431 11450
rect 18431 11398 18443 11450
rect 18443 11398 18457 11450
rect 18481 11398 18495 11450
rect 18495 11398 18507 11450
rect 18507 11398 18537 11450
rect 18561 11398 18571 11450
rect 18571 11398 18617 11450
rect 18321 11396 18377 11398
rect 18401 11396 18457 11398
rect 18481 11396 18537 11398
rect 18561 11396 18617 11398
rect 18321 10362 18377 10364
rect 18401 10362 18457 10364
rect 18481 10362 18537 10364
rect 18561 10362 18617 10364
rect 18321 10310 18367 10362
rect 18367 10310 18377 10362
rect 18401 10310 18431 10362
rect 18431 10310 18443 10362
rect 18443 10310 18457 10362
rect 18481 10310 18495 10362
rect 18495 10310 18507 10362
rect 18507 10310 18537 10362
rect 18561 10310 18571 10362
rect 18571 10310 18617 10362
rect 18321 10308 18377 10310
rect 18401 10308 18457 10310
rect 18481 10308 18537 10310
rect 18561 10308 18617 10310
rect 17774 9424 17830 9480
rect 17774 9288 17830 9344
rect 17130 4140 17186 4176
rect 17130 4120 17132 4140
rect 17132 4120 17184 4140
rect 17184 4120 17186 4140
rect 17774 7828 17776 7848
rect 17776 7828 17828 7848
rect 17828 7828 17830 7848
rect 17774 7792 17830 7828
rect 17866 7248 17922 7304
rect 18321 9274 18377 9276
rect 18401 9274 18457 9276
rect 18481 9274 18537 9276
rect 18561 9274 18617 9276
rect 18321 9222 18367 9274
rect 18367 9222 18377 9274
rect 18401 9222 18431 9274
rect 18431 9222 18443 9274
rect 18443 9222 18457 9274
rect 18481 9222 18495 9274
rect 18495 9222 18507 9274
rect 18507 9222 18537 9274
rect 18561 9222 18571 9274
rect 18571 9222 18617 9274
rect 18321 9220 18377 9222
rect 18401 9220 18457 9222
rect 18481 9220 18537 9222
rect 18561 9220 18617 9222
rect 18981 10906 19037 10908
rect 19061 10906 19117 10908
rect 19141 10906 19197 10908
rect 19221 10906 19277 10908
rect 18981 10854 19027 10906
rect 19027 10854 19037 10906
rect 19061 10854 19091 10906
rect 19091 10854 19103 10906
rect 19103 10854 19117 10906
rect 19141 10854 19155 10906
rect 19155 10854 19167 10906
rect 19167 10854 19197 10906
rect 19221 10854 19231 10906
rect 19231 10854 19277 10906
rect 18981 10852 19037 10854
rect 19061 10852 19117 10854
rect 19141 10852 19197 10854
rect 19221 10852 19277 10854
rect 18981 9818 19037 9820
rect 19061 9818 19117 9820
rect 19141 9818 19197 9820
rect 19221 9818 19277 9820
rect 18981 9766 19027 9818
rect 19027 9766 19037 9818
rect 19061 9766 19091 9818
rect 19091 9766 19103 9818
rect 19103 9766 19117 9818
rect 19141 9766 19155 9818
rect 19155 9766 19167 9818
rect 19167 9766 19197 9818
rect 19221 9766 19231 9818
rect 19231 9766 19277 9818
rect 18981 9764 19037 9766
rect 19061 9764 19117 9766
rect 19141 9764 19197 9766
rect 19221 9764 19277 9766
rect 18321 8186 18377 8188
rect 18401 8186 18457 8188
rect 18481 8186 18537 8188
rect 18561 8186 18617 8188
rect 18321 8134 18367 8186
rect 18367 8134 18377 8186
rect 18401 8134 18431 8186
rect 18431 8134 18443 8186
rect 18443 8134 18457 8186
rect 18481 8134 18495 8186
rect 18495 8134 18507 8186
rect 18507 8134 18537 8186
rect 18561 8134 18571 8186
rect 18571 8134 18617 8186
rect 18321 8132 18377 8134
rect 18401 8132 18457 8134
rect 18481 8132 18537 8134
rect 18561 8132 18617 8134
rect 18694 7828 18696 7848
rect 18696 7828 18748 7848
rect 18748 7828 18750 7848
rect 18694 7792 18750 7828
rect 18321 7098 18377 7100
rect 18401 7098 18457 7100
rect 18481 7098 18537 7100
rect 18561 7098 18617 7100
rect 18321 7046 18367 7098
rect 18367 7046 18377 7098
rect 18401 7046 18431 7098
rect 18431 7046 18443 7098
rect 18443 7046 18457 7098
rect 18481 7046 18495 7098
rect 18495 7046 18507 7098
rect 18507 7046 18537 7098
rect 18561 7046 18571 7098
rect 18571 7046 18617 7098
rect 18321 7044 18377 7046
rect 18401 7044 18457 7046
rect 18481 7044 18537 7046
rect 18561 7044 18617 7046
rect 18878 9036 18934 9072
rect 18878 9016 18880 9036
rect 18880 9016 18932 9036
rect 18932 9016 18934 9036
rect 18981 8730 19037 8732
rect 19061 8730 19117 8732
rect 19141 8730 19197 8732
rect 19221 8730 19277 8732
rect 18981 8678 19027 8730
rect 19027 8678 19037 8730
rect 19061 8678 19091 8730
rect 19091 8678 19103 8730
rect 19103 8678 19117 8730
rect 19141 8678 19155 8730
rect 19155 8678 19167 8730
rect 19167 8678 19197 8730
rect 19221 8678 19231 8730
rect 19231 8678 19277 8730
rect 18981 8676 19037 8678
rect 19061 8676 19117 8678
rect 19141 8676 19197 8678
rect 19221 8676 19277 8678
rect 18981 7642 19037 7644
rect 19061 7642 19117 7644
rect 19141 7642 19197 7644
rect 19221 7642 19277 7644
rect 18981 7590 19027 7642
rect 19027 7590 19037 7642
rect 19061 7590 19091 7642
rect 19091 7590 19103 7642
rect 19103 7590 19117 7642
rect 19141 7590 19155 7642
rect 19155 7590 19167 7642
rect 19167 7590 19197 7642
rect 19221 7590 19231 7642
rect 19231 7590 19277 7642
rect 18981 7588 19037 7590
rect 19061 7588 19117 7590
rect 19141 7588 19197 7590
rect 19221 7588 19277 7590
rect 25267 27770 25323 27772
rect 25347 27770 25403 27772
rect 25427 27770 25483 27772
rect 25507 27770 25563 27772
rect 25267 27718 25313 27770
rect 25313 27718 25323 27770
rect 25347 27718 25377 27770
rect 25377 27718 25389 27770
rect 25389 27718 25403 27770
rect 25427 27718 25441 27770
rect 25441 27718 25453 27770
rect 25453 27718 25483 27770
rect 25507 27718 25517 27770
rect 25517 27718 25563 27770
rect 25267 27716 25323 27718
rect 25347 27716 25403 27718
rect 25427 27716 25483 27718
rect 25507 27716 25563 27718
rect 25927 27226 25983 27228
rect 26007 27226 26063 27228
rect 26087 27226 26143 27228
rect 26167 27226 26223 27228
rect 25927 27174 25973 27226
rect 25973 27174 25983 27226
rect 26007 27174 26037 27226
rect 26037 27174 26049 27226
rect 26049 27174 26063 27226
rect 26087 27174 26101 27226
rect 26101 27174 26113 27226
rect 26113 27174 26143 27226
rect 26167 27174 26177 27226
rect 26177 27174 26223 27226
rect 25927 27172 25983 27174
rect 26007 27172 26063 27174
rect 26087 27172 26143 27174
rect 26167 27172 26223 27174
rect 25267 26682 25323 26684
rect 25347 26682 25403 26684
rect 25427 26682 25483 26684
rect 25507 26682 25563 26684
rect 25267 26630 25313 26682
rect 25313 26630 25323 26682
rect 25347 26630 25377 26682
rect 25377 26630 25389 26682
rect 25389 26630 25403 26682
rect 25427 26630 25441 26682
rect 25441 26630 25453 26682
rect 25453 26630 25483 26682
rect 25507 26630 25517 26682
rect 25517 26630 25563 26682
rect 25267 26628 25323 26630
rect 25347 26628 25403 26630
rect 25427 26628 25483 26630
rect 25507 26628 25563 26630
rect 25927 26138 25983 26140
rect 26007 26138 26063 26140
rect 26087 26138 26143 26140
rect 26167 26138 26223 26140
rect 25927 26086 25973 26138
rect 25973 26086 25983 26138
rect 26007 26086 26037 26138
rect 26037 26086 26049 26138
rect 26049 26086 26063 26138
rect 26087 26086 26101 26138
rect 26101 26086 26113 26138
rect 26113 26086 26143 26138
rect 26167 26086 26177 26138
rect 26177 26086 26223 26138
rect 25927 26084 25983 26086
rect 26007 26084 26063 26086
rect 26087 26084 26143 26086
rect 26167 26084 26223 26086
rect 25267 25594 25323 25596
rect 25347 25594 25403 25596
rect 25427 25594 25483 25596
rect 25507 25594 25563 25596
rect 25267 25542 25313 25594
rect 25313 25542 25323 25594
rect 25347 25542 25377 25594
rect 25377 25542 25389 25594
rect 25389 25542 25403 25594
rect 25427 25542 25441 25594
rect 25441 25542 25453 25594
rect 25453 25542 25483 25594
rect 25507 25542 25517 25594
rect 25517 25542 25563 25594
rect 25267 25540 25323 25542
rect 25347 25540 25403 25542
rect 25427 25540 25483 25542
rect 25507 25540 25563 25542
rect 28538 25236 28540 25256
rect 28540 25236 28592 25256
rect 28592 25236 28594 25256
rect 25927 25050 25983 25052
rect 26007 25050 26063 25052
rect 26087 25050 26143 25052
rect 26167 25050 26223 25052
rect 25927 24998 25973 25050
rect 25973 24998 25983 25050
rect 26007 24998 26037 25050
rect 26037 24998 26049 25050
rect 26049 24998 26063 25050
rect 26087 24998 26101 25050
rect 26101 24998 26113 25050
rect 26113 24998 26143 25050
rect 26167 24998 26177 25050
rect 26177 24998 26223 25050
rect 25927 24996 25983 24998
rect 26007 24996 26063 24998
rect 26087 24996 26143 24998
rect 26167 24996 26223 24998
rect 25267 24506 25323 24508
rect 25347 24506 25403 24508
rect 25427 24506 25483 24508
rect 25507 24506 25563 24508
rect 25267 24454 25313 24506
rect 25313 24454 25323 24506
rect 25347 24454 25377 24506
rect 25377 24454 25389 24506
rect 25389 24454 25403 24506
rect 25427 24454 25441 24506
rect 25441 24454 25453 24506
rect 25453 24454 25483 24506
rect 25507 24454 25517 24506
rect 25517 24454 25563 24506
rect 25267 24452 25323 24454
rect 25347 24452 25403 24454
rect 25427 24452 25483 24454
rect 25507 24452 25563 24454
rect 25927 23962 25983 23964
rect 26007 23962 26063 23964
rect 26087 23962 26143 23964
rect 26167 23962 26223 23964
rect 25927 23910 25973 23962
rect 25973 23910 25983 23962
rect 26007 23910 26037 23962
rect 26037 23910 26049 23962
rect 26049 23910 26063 23962
rect 26087 23910 26101 23962
rect 26101 23910 26113 23962
rect 26113 23910 26143 23962
rect 26167 23910 26177 23962
rect 26177 23910 26223 23962
rect 25927 23908 25983 23910
rect 26007 23908 26063 23910
rect 26087 23908 26143 23910
rect 26167 23908 26223 23910
rect 25267 23418 25323 23420
rect 25347 23418 25403 23420
rect 25427 23418 25483 23420
rect 25507 23418 25563 23420
rect 25267 23366 25313 23418
rect 25313 23366 25323 23418
rect 25347 23366 25377 23418
rect 25377 23366 25389 23418
rect 25389 23366 25403 23418
rect 25427 23366 25441 23418
rect 25441 23366 25453 23418
rect 25453 23366 25483 23418
rect 25507 23366 25517 23418
rect 25517 23366 25563 23418
rect 25267 23364 25323 23366
rect 25347 23364 25403 23366
rect 25427 23364 25483 23366
rect 25507 23364 25563 23366
rect 25927 22874 25983 22876
rect 26007 22874 26063 22876
rect 26087 22874 26143 22876
rect 26167 22874 26223 22876
rect 25927 22822 25973 22874
rect 25973 22822 25983 22874
rect 26007 22822 26037 22874
rect 26037 22822 26049 22874
rect 26049 22822 26063 22874
rect 26087 22822 26101 22874
rect 26101 22822 26113 22874
rect 26113 22822 26143 22874
rect 26167 22822 26177 22874
rect 26177 22822 26223 22874
rect 25927 22820 25983 22822
rect 26007 22820 26063 22822
rect 26087 22820 26143 22822
rect 26167 22820 26223 22822
rect 25267 22330 25323 22332
rect 25347 22330 25403 22332
rect 25427 22330 25483 22332
rect 25507 22330 25563 22332
rect 25267 22278 25313 22330
rect 25313 22278 25323 22330
rect 25347 22278 25377 22330
rect 25377 22278 25389 22330
rect 25389 22278 25403 22330
rect 25427 22278 25441 22330
rect 25441 22278 25453 22330
rect 25453 22278 25483 22330
rect 25507 22278 25517 22330
rect 25517 22278 25563 22330
rect 25267 22276 25323 22278
rect 25347 22276 25403 22278
rect 25427 22276 25483 22278
rect 25507 22276 25563 22278
rect 25927 21786 25983 21788
rect 26007 21786 26063 21788
rect 26087 21786 26143 21788
rect 26167 21786 26223 21788
rect 25927 21734 25973 21786
rect 25973 21734 25983 21786
rect 26007 21734 26037 21786
rect 26037 21734 26049 21786
rect 26049 21734 26063 21786
rect 26087 21734 26101 21786
rect 26101 21734 26113 21786
rect 26113 21734 26143 21786
rect 26167 21734 26177 21786
rect 26177 21734 26223 21786
rect 25927 21732 25983 21734
rect 26007 21732 26063 21734
rect 26087 21732 26143 21734
rect 26167 21732 26223 21734
rect 25267 21242 25323 21244
rect 25347 21242 25403 21244
rect 25427 21242 25483 21244
rect 25507 21242 25563 21244
rect 25267 21190 25313 21242
rect 25313 21190 25323 21242
rect 25347 21190 25377 21242
rect 25377 21190 25389 21242
rect 25389 21190 25403 21242
rect 25427 21190 25441 21242
rect 25441 21190 25453 21242
rect 25453 21190 25483 21242
rect 25507 21190 25517 21242
rect 25517 21190 25563 21242
rect 25267 21188 25323 21190
rect 25347 21188 25403 21190
rect 25427 21188 25483 21190
rect 25507 21188 25563 21190
rect 25927 20698 25983 20700
rect 26007 20698 26063 20700
rect 26087 20698 26143 20700
rect 26167 20698 26223 20700
rect 25927 20646 25973 20698
rect 25973 20646 25983 20698
rect 26007 20646 26037 20698
rect 26037 20646 26049 20698
rect 26049 20646 26063 20698
rect 26087 20646 26101 20698
rect 26101 20646 26113 20698
rect 26113 20646 26143 20698
rect 26167 20646 26177 20698
rect 26177 20646 26223 20698
rect 25927 20644 25983 20646
rect 26007 20644 26063 20646
rect 26087 20644 26143 20646
rect 26167 20644 26223 20646
rect 25267 20154 25323 20156
rect 25347 20154 25403 20156
rect 25427 20154 25483 20156
rect 25507 20154 25563 20156
rect 25267 20102 25313 20154
rect 25313 20102 25323 20154
rect 25347 20102 25377 20154
rect 25377 20102 25389 20154
rect 25389 20102 25403 20154
rect 25427 20102 25441 20154
rect 25441 20102 25453 20154
rect 25453 20102 25483 20154
rect 25507 20102 25517 20154
rect 25517 20102 25563 20154
rect 25267 20100 25323 20102
rect 25347 20100 25403 20102
rect 25427 20100 25483 20102
rect 25507 20100 25563 20102
rect 25927 19610 25983 19612
rect 26007 19610 26063 19612
rect 26087 19610 26143 19612
rect 26167 19610 26223 19612
rect 25927 19558 25973 19610
rect 25973 19558 25983 19610
rect 26007 19558 26037 19610
rect 26037 19558 26049 19610
rect 26049 19558 26063 19610
rect 26087 19558 26101 19610
rect 26101 19558 26113 19610
rect 26113 19558 26143 19610
rect 26167 19558 26177 19610
rect 26177 19558 26223 19610
rect 25927 19556 25983 19558
rect 26007 19556 26063 19558
rect 26087 19556 26143 19558
rect 26167 19556 26223 19558
rect 25267 19066 25323 19068
rect 25347 19066 25403 19068
rect 25427 19066 25483 19068
rect 25507 19066 25563 19068
rect 25267 19014 25313 19066
rect 25313 19014 25323 19066
rect 25347 19014 25377 19066
rect 25377 19014 25389 19066
rect 25389 19014 25403 19066
rect 25427 19014 25441 19066
rect 25441 19014 25453 19066
rect 25453 19014 25483 19066
rect 25507 19014 25517 19066
rect 25517 19014 25563 19066
rect 25267 19012 25323 19014
rect 25347 19012 25403 19014
rect 25427 19012 25483 19014
rect 25507 19012 25563 19014
rect 25927 18522 25983 18524
rect 26007 18522 26063 18524
rect 26087 18522 26143 18524
rect 26167 18522 26223 18524
rect 25927 18470 25973 18522
rect 25973 18470 25983 18522
rect 26007 18470 26037 18522
rect 26037 18470 26049 18522
rect 26049 18470 26063 18522
rect 26087 18470 26101 18522
rect 26101 18470 26113 18522
rect 26113 18470 26143 18522
rect 26167 18470 26177 18522
rect 26177 18470 26223 18522
rect 25927 18468 25983 18470
rect 26007 18468 26063 18470
rect 26087 18468 26143 18470
rect 26167 18468 26223 18470
rect 25267 17978 25323 17980
rect 25347 17978 25403 17980
rect 25427 17978 25483 17980
rect 25507 17978 25563 17980
rect 25267 17926 25313 17978
rect 25313 17926 25323 17978
rect 25347 17926 25377 17978
rect 25377 17926 25389 17978
rect 25389 17926 25403 17978
rect 25427 17926 25441 17978
rect 25441 17926 25453 17978
rect 25453 17926 25483 17978
rect 25507 17926 25517 17978
rect 25517 17926 25563 17978
rect 25267 17924 25323 17926
rect 25347 17924 25403 17926
rect 25427 17924 25483 17926
rect 25507 17924 25563 17926
rect 25927 17434 25983 17436
rect 26007 17434 26063 17436
rect 26087 17434 26143 17436
rect 26167 17434 26223 17436
rect 25927 17382 25973 17434
rect 25973 17382 25983 17434
rect 26007 17382 26037 17434
rect 26037 17382 26049 17434
rect 26049 17382 26063 17434
rect 26087 17382 26101 17434
rect 26101 17382 26113 17434
rect 26113 17382 26143 17434
rect 26167 17382 26177 17434
rect 26177 17382 26223 17434
rect 25927 17380 25983 17382
rect 26007 17380 26063 17382
rect 26087 17380 26143 17382
rect 26167 17380 26223 17382
rect 25267 16890 25323 16892
rect 25347 16890 25403 16892
rect 25427 16890 25483 16892
rect 25507 16890 25563 16892
rect 25267 16838 25313 16890
rect 25313 16838 25323 16890
rect 25347 16838 25377 16890
rect 25377 16838 25389 16890
rect 25389 16838 25403 16890
rect 25427 16838 25441 16890
rect 25441 16838 25453 16890
rect 25453 16838 25483 16890
rect 25507 16838 25517 16890
rect 25517 16838 25563 16890
rect 25267 16836 25323 16838
rect 25347 16836 25403 16838
rect 25427 16836 25483 16838
rect 25507 16836 25563 16838
rect 25927 16346 25983 16348
rect 26007 16346 26063 16348
rect 26087 16346 26143 16348
rect 26167 16346 26223 16348
rect 25927 16294 25973 16346
rect 25973 16294 25983 16346
rect 26007 16294 26037 16346
rect 26037 16294 26049 16346
rect 26049 16294 26063 16346
rect 26087 16294 26101 16346
rect 26101 16294 26113 16346
rect 26113 16294 26143 16346
rect 26167 16294 26177 16346
rect 26177 16294 26223 16346
rect 25927 16292 25983 16294
rect 26007 16292 26063 16294
rect 26087 16292 26143 16294
rect 26167 16292 26223 16294
rect 25267 15802 25323 15804
rect 25347 15802 25403 15804
rect 25427 15802 25483 15804
rect 25507 15802 25563 15804
rect 25267 15750 25313 15802
rect 25313 15750 25323 15802
rect 25347 15750 25377 15802
rect 25377 15750 25389 15802
rect 25389 15750 25403 15802
rect 25427 15750 25441 15802
rect 25441 15750 25453 15802
rect 25453 15750 25483 15802
rect 25507 15750 25517 15802
rect 25517 15750 25563 15802
rect 25267 15748 25323 15750
rect 25347 15748 25403 15750
rect 25427 15748 25483 15750
rect 25507 15748 25563 15750
rect 25927 15258 25983 15260
rect 26007 15258 26063 15260
rect 26087 15258 26143 15260
rect 26167 15258 26223 15260
rect 25927 15206 25973 15258
rect 25973 15206 25983 15258
rect 26007 15206 26037 15258
rect 26037 15206 26049 15258
rect 26049 15206 26063 15258
rect 26087 15206 26101 15258
rect 26101 15206 26113 15258
rect 26113 15206 26143 15258
rect 26167 15206 26177 15258
rect 26177 15206 26223 15258
rect 25927 15204 25983 15206
rect 26007 15204 26063 15206
rect 26087 15204 26143 15206
rect 26167 15204 26223 15206
rect 25267 14714 25323 14716
rect 25347 14714 25403 14716
rect 25427 14714 25483 14716
rect 25507 14714 25563 14716
rect 25267 14662 25313 14714
rect 25313 14662 25323 14714
rect 25347 14662 25377 14714
rect 25377 14662 25389 14714
rect 25389 14662 25403 14714
rect 25427 14662 25441 14714
rect 25441 14662 25453 14714
rect 25453 14662 25483 14714
rect 25507 14662 25517 14714
rect 25517 14662 25563 14714
rect 25267 14660 25323 14662
rect 25347 14660 25403 14662
rect 25427 14660 25483 14662
rect 25507 14660 25563 14662
rect 25927 14170 25983 14172
rect 26007 14170 26063 14172
rect 26087 14170 26143 14172
rect 26167 14170 26223 14172
rect 25927 14118 25973 14170
rect 25973 14118 25983 14170
rect 26007 14118 26037 14170
rect 26037 14118 26049 14170
rect 26049 14118 26063 14170
rect 26087 14118 26101 14170
rect 26101 14118 26113 14170
rect 26113 14118 26143 14170
rect 26167 14118 26177 14170
rect 26177 14118 26223 14170
rect 25927 14116 25983 14118
rect 26007 14116 26063 14118
rect 26087 14116 26143 14118
rect 26167 14116 26223 14118
rect 25267 13626 25323 13628
rect 25347 13626 25403 13628
rect 25427 13626 25483 13628
rect 25507 13626 25563 13628
rect 25267 13574 25313 13626
rect 25313 13574 25323 13626
rect 25347 13574 25377 13626
rect 25377 13574 25389 13626
rect 25389 13574 25403 13626
rect 25427 13574 25441 13626
rect 25441 13574 25453 13626
rect 25453 13574 25483 13626
rect 25507 13574 25517 13626
rect 25517 13574 25563 13626
rect 25267 13572 25323 13574
rect 25347 13572 25403 13574
rect 25427 13572 25483 13574
rect 25507 13572 25563 13574
rect 25927 13082 25983 13084
rect 26007 13082 26063 13084
rect 26087 13082 26143 13084
rect 26167 13082 26223 13084
rect 25927 13030 25973 13082
rect 25973 13030 25983 13082
rect 26007 13030 26037 13082
rect 26037 13030 26049 13082
rect 26049 13030 26063 13082
rect 26087 13030 26101 13082
rect 26101 13030 26113 13082
rect 26113 13030 26143 13082
rect 26167 13030 26177 13082
rect 26177 13030 26223 13082
rect 25927 13028 25983 13030
rect 26007 13028 26063 13030
rect 26087 13028 26143 13030
rect 26167 13028 26223 13030
rect 28538 25200 28594 25236
rect 25267 12538 25323 12540
rect 25347 12538 25403 12540
rect 25427 12538 25483 12540
rect 25507 12538 25563 12540
rect 25267 12486 25313 12538
rect 25313 12486 25323 12538
rect 25347 12486 25377 12538
rect 25377 12486 25389 12538
rect 25389 12486 25403 12538
rect 25427 12486 25441 12538
rect 25441 12486 25453 12538
rect 25453 12486 25483 12538
rect 25507 12486 25517 12538
rect 25517 12486 25563 12538
rect 25267 12484 25323 12486
rect 25347 12484 25403 12486
rect 25427 12484 25483 12486
rect 25507 12484 25563 12486
rect 25927 11994 25983 11996
rect 26007 11994 26063 11996
rect 26087 11994 26143 11996
rect 26167 11994 26223 11996
rect 25927 11942 25973 11994
rect 25973 11942 25983 11994
rect 26007 11942 26037 11994
rect 26037 11942 26049 11994
rect 26049 11942 26063 11994
rect 26087 11942 26101 11994
rect 26101 11942 26113 11994
rect 26113 11942 26143 11994
rect 26167 11942 26177 11994
rect 26177 11942 26223 11994
rect 25927 11940 25983 11942
rect 26007 11940 26063 11942
rect 26087 11940 26143 11942
rect 26167 11940 26223 11942
rect 5089 2202 5145 2204
rect 5169 2202 5225 2204
rect 5249 2202 5305 2204
rect 5329 2202 5385 2204
rect 5089 2150 5135 2202
rect 5135 2150 5145 2202
rect 5169 2150 5199 2202
rect 5199 2150 5211 2202
rect 5211 2150 5225 2202
rect 5249 2150 5263 2202
rect 5263 2150 5275 2202
rect 5275 2150 5305 2202
rect 5329 2150 5339 2202
rect 5339 2150 5385 2202
rect 5089 2148 5145 2150
rect 5169 2148 5225 2150
rect 5249 2148 5305 2150
rect 5329 2148 5385 2150
rect 18321 6010 18377 6012
rect 18401 6010 18457 6012
rect 18481 6010 18537 6012
rect 18561 6010 18617 6012
rect 18321 5958 18367 6010
rect 18367 5958 18377 6010
rect 18401 5958 18431 6010
rect 18431 5958 18443 6010
rect 18443 5958 18457 6010
rect 18481 5958 18495 6010
rect 18495 5958 18507 6010
rect 18507 5958 18537 6010
rect 18561 5958 18571 6010
rect 18571 5958 18617 6010
rect 18321 5956 18377 5958
rect 18401 5956 18457 5958
rect 18481 5956 18537 5958
rect 18561 5956 18617 5958
rect 18321 4922 18377 4924
rect 18401 4922 18457 4924
rect 18481 4922 18537 4924
rect 18561 4922 18617 4924
rect 18321 4870 18367 4922
rect 18367 4870 18377 4922
rect 18401 4870 18431 4922
rect 18431 4870 18443 4922
rect 18443 4870 18457 4922
rect 18481 4870 18495 4922
rect 18495 4870 18507 4922
rect 18507 4870 18537 4922
rect 18561 4870 18571 4922
rect 18571 4870 18617 4922
rect 18321 4868 18377 4870
rect 18401 4868 18457 4870
rect 18481 4868 18537 4870
rect 18561 4868 18617 4870
rect 18981 6554 19037 6556
rect 19061 6554 19117 6556
rect 19141 6554 19197 6556
rect 19221 6554 19277 6556
rect 18981 6502 19027 6554
rect 19027 6502 19037 6554
rect 19061 6502 19091 6554
rect 19091 6502 19103 6554
rect 19103 6502 19117 6554
rect 19141 6502 19155 6554
rect 19155 6502 19167 6554
rect 19167 6502 19197 6554
rect 19221 6502 19231 6554
rect 19231 6502 19277 6554
rect 18981 6500 19037 6502
rect 19061 6500 19117 6502
rect 19141 6500 19197 6502
rect 19221 6500 19277 6502
rect 20810 7248 20866 7304
rect 18981 5466 19037 5468
rect 19061 5466 19117 5468
rect 19141 5466 19197 5468
rect 19221 5466 19277 5468
rect 18981 5414 19027 5466
rect 19027 5414 19037 5466
rect 19061 5414 19091 5466
rect 19091 5414 19103 5466
rect 19103 5414 19117 5466
rect 19141 5414 19155 5466
rect 19155 5414 19167 5466
rect 19167 5414 19197 5466
rect 19221 5414 19231 5466
rect 19231 5414 19277 5466
rect 18981 5412 19037 5414
rect 19061 5412 19117 5414
rect 19141 5412 19197 5414
rect 19221 5412 19277 5414
rect 18321 3834 18377 3836
rect 18401 3834 18457 3836
rect 18481 3834 18537 3836
rect 18561 3834 18617 3836
rect 18321 3782 18367 3834
rect 18367 3782 18377 3834
rect 18401 3782 18431 3834
rect 18431 3782 18443 3834
rect 18443 3782 18457 3834
rect 18481 3782 18495 3834
rect 18495 3782 18507 3834
rect 18507 3782 18537 3834
rect 18561 3782 18571 3834
rect 18571 3782 18617 3834
rect 18321 3780 18377 3782
rect 18401 3780 18457 3782
rect 18481 3780 18537 3782
rect 18561 3780 18617 3782
rect 18321 2746 18377 2748
rect 18401 2746 18457 2748
rect 18481 2746 18537 2748
rect 18561 2746 18617 2748
rect 18321 2694 18367 2746
rect 18367 2694 18377 2746
rect 18401 2694 18431 2746
rect 18431 2694 18443 2746
rect 18443 2694 18457 2746
rect 18481 2694 18495 2746
rect 18495 2694 18507 2746
rect 18507 2694 18537 2746
rect 18561 2694 18571 2746
rect 18571 2694 18617 2746
rect 18321 2692 18377 2694
rect 18401 2692 18457 2694
rect 18481 2692 18537 2694
rect 18561 2692 18617 2694
rect 12035 2202 12091 2204
rect 12115 2202 12171 2204
rect 12195 2202 12251 2204
rect 12275 2202 12331 2204
rect 12035 2150 12081 2202
rect 12081 2150 12091 2202
rect 12115 2150 12145 2202
rect 12145 2150 12157 2202
rect 12157 2150 12171 2202
rect 12195 2150 12209 2202
rect 12209 2150 12221 2202
rect 12221 2150 12251 2202
rect 12275 2150 12285 2202
rect 12285 2150 12331 2202
rect 12035 2148 12091 2150
rect 12115 2148 12171 2150
rect 12195 2148 12251 2150
rect 12275 2148 12331 2150
rect 18981 4378 19037 4380
rect 19061 4378 19117 4380
rect 19141 4378 19197 4380
rect 19221 4378 19277 4380
rect 18981 4326 19027 4378
rect 19027 4326 19037 4378
rect 19061 4326 19091 4378
rect 19091 4326 19103 4378
rect 19103 4326 19117 4378
rect 19141 4326 19155 4378
rect 19155 4326 19167 4378
rect 19167 4326 19197 4378
rect 19221 4326 19231 4378
rect 19231 4326 19277 4378
rect 18981 4324 19037 4326
rect 19061 4324 19117 4326
rect 19141 4324 19197 4326
rect 19221 4324 19277 4326
rect 18970 4140 19026 4176
rect 18970 4120 18972 4140
rect 18972 4120 19024 4140
rect 19024 4120 19026 4140
rect 18981 3290 19037 3292
rect 19061 3290 19117 3292
rect 19141 3290 19197 3292
rect 19221 3290 19277 3292
rect 18981 3238 19027 3290
rect 19027 3238 19037 3290
rect 19061 3238 19091 3290
rect 19091 3238 19103 3290
rect 19103 3238 19117 3290
rect 19141 3238 19155 3290
rect 19155 3238 19167 3290
rect 19167 3238 19197 3290
rect 19221 3238 19231 3290
rect 19231 3238 19277 3290
rect 18981 3236 19037 3238
rect 19061 3236 19117 3238
rect 19141 3236 19197 3238
rect 19221 3236 19277 3238
rect 25267 11450 25323 11452
rect 25347 11450 25403 11452
rect 25427 11450 25483 11452
rect 25507 11450 25563 11452
rect 25267 11398 25313 11450
rect 25313 11398 25323 11450
rect 25347 11398 25377 11450
rect 25377 11398 25389 11450
rect 25389 11398 25403 11450
rect 25427 11398 25441 11450
rect 25441 11398 25453 11450
rect 25453 11398 25483 11450
rect 25507 11398 25517 11450
rect 25517 11398 25563 11450
rect 25267 11396 25323 11398
rect 25347 11396 25403 11398
rect 25427 11396 25483 11398
rect 25507 11396 25563 11398
rect 25927 10906 25983 10908
rect 26007 10906 26063 10908
rect 26087 10906 26143 10908
rect 26167 10906 26223 10908
rect 25927 10854 25973 10906
rect 25973 10854 25983 10906
rect 26007 10854 26037 10906
rect 26037 10854 26049 10906
rect 26049 10854 26063 10906
rect 26087 10854 26101 10906
rect 26101 10854 26113 10906
rect 26113 10854 26143 10906
rect 26167 10854 26177 10906
rect 26177 10854 26223 10906
rect 25927 10852 25983 10854
rect 26007 10852 26063 10854
rect 26087 10852 26143 10854
rect 26167 10852 26223 10854
rect 21822 8200 21878 8256
rect 21914 7248 21970 7304
rect 25267 10362 25323 10364
rect 25347 10362 25403 10364
rect 25427 10362 25483 10364
rect 25507 10362 25563 10364
rect 25267 10310 25313 10362
rect 25313 10310 25323 10362
rect 25347 10310 25377 10362
rect 25377 10310 25389 10362
rect 25389 10310 25403 10362
rect 25427 10310 25441 10362
rect 25441 10310 25453 10362
rect 25453 10310 25483 10362
rect 25507 10310 25517 10362
rect 25517 10310 25563 10362
rect 25267 10308 25323 10310
rect 25347 10308 25403 10310
rect 25427 10308 25483 10310
rect 25507 10308 25563 10310
rect 25927 9818 25983 9820
rect 26007 9818 26063 9820
rect 26087 9818 26143 9820
rect 26167 9818 26223 9820
rect 25927 9766 25973 9818
rect 25973 9766 25983 9818
rect 26007 9766 26037 9818
rect 26037 9766 26049 9818
rect 26049 9766 26063 9818
rect 26087 9766 26101 9818
rect 26101 9766 26113 9818
rect 26113 9766 26143 9818
rect 26167 9766 26177 9818
rect 26177 9766 26223 9818
rect 25927 9764 25983 9766
rect 26007 9764 26063 9766
rect 26087 9764 26143 9766
rect 26167 9764 26223 9766
rect 25267 9274 25323 9276
rect 25347 9274 25403 9276
rect 25427 9274 25483 9276
rect 25507 9274 25563 9276
rect 25267 9222 25313 9274
rect 25313 9222 25323 9274
rect 25347 9222 25377 9274
rect 25377 9222 25389 9274
rect 25389 9222 25403 9274
rect 25427 9222 25441 9274
rect 25441 9222 25453 9274
rect 25453 9222 25483 9274
rect 25507 9222 25517 9274
rect 25517 9222 25563 9274
rect 25267 9220 25323 9222
rect 25347 9220 25403 9222
rect 25427 9220 25483 9222
rect 25507 9220 25563 9222
rect 25927 8730 25983 8732
rect 26007 8730 26063 8732
rect 26087 8730 26143 8732
rect 26167 8730 26223 8732
rect 25927 8678 25973 8730
rect 25973 8678 25983 8730
rect 26007 8678 26037 8730
rect 26037 8678 26049 8730
rect 26049 8678 26063 8730
rect 26087 8678 26101 8730
rect 26101 8678 26113 8730
rect 26113 8678 26143 8730
rect 26167 8678 26177 8730
rect 26177 8678 26223 8730
rect 25927 8676 25983 8678
rect 26007 8676 26063 8678
rect 26087 8676 26143 8678
rect 26167 8676 26223 8678
rect 25267 8186 25323 8188
rect 25347 8186 25403 8188
rect 25427 8186 25483 8188
rect 25507 8186 25563 8188
rect 25267 8134 25313 8186
rect 25313 8134 25323 8186
rect 25347 8134 25377 8186
rect 25377 8134 25389 8186
rect 25389 8134 25403 8186
rect 25427 8134 25441 8186
rect 25441 8134 25453 8186
rect 25453 8134 25483 8186
rect 25507 8134 25517 8186
rect 25517 8134 25563 8186
rect 25267 8132 25323 8134
rect 25347 8132 25403 8134
rect 25427 8132 25483 8134
rect 25507 8132 25563 8134
rect 22926 7248 22982 7304
rect 25927 7642 25983 7644
rect 26007 7642 26063 7644
rect 26087 7642 26143 7644
rect 26167 7642 26223 7644
rect 25927 7590 25973 7642
rect 25973 7590 25983 7642
rect 26007 7590 26037 7642
rect 26037 7590 26049 7642
rect 26049 7590 26063 7642
rect 26087 7590 26101 7642
rect 26101 7590 26113 7642
rect 26113 7590 26143 7642
rect 26167 7590 26177 7642
rect 26177 7590 26223 7642
rect 25927 7588 25983 7590
rect 26007 7588 26063 7590
rect 26087 7588 26143 7590
rect 26167 7588 26223 7590
rect 25267 7098 25323 7100
rect 25347 7098 25403 7100
rect 25427 7098 25483 7100
rect 25507 7098 25563 7100
rect 25267 7046 25313 7098
rect 25313 7046 25323 7098
rect 25347 7046 25377 7098
rect 25377 7046 25389 7098
rect 25389 7046 25403 7098
rect 25427 7046 25441 7098
rect 25441 7046 25453 7098
rect 25453 7046 25483 7098
rect 25507 7046 25517 7098
rect 25517 7046 25563 7098
rect 25267 7044 25323 7046
rect 25347 7044 25403 7046
rect 25427 7044 25483 7046
rect 25507 7044 25563 7046
rect 25267 6010 25323 6012
rect 25347 6010 25403 6012
rect 25427 6010 25483 6012
rect 25507 6010 25563 6012
rect 25267 5958 25313 6010
rect 25313 5958 25323 6010
rect 25347 5958 25377 6010
rect 25377 5958 25389 6010
rect 25389 5958 25403 6010
rect 25427 5958 25441 6010
rect 25441 5958 25453 6010
rect 25453 5958 25483 6010
rect 25507 5958 25517 6010
rect 25517 5958 25563 6010
rect 25267 5956 25323 5958
rect 25347 5956 25403 5958
rect 25427 5956 25483 5958
rect 25507 5956 25563 5958
rect 25927 6554 25983 6556
rect 26007 6554 26063 6556
rect 26087 6554 26143 6556
rect 26167 6554 26223 6556
rect 25927 6502 25973 6554
rect 25973 6502 25983 6554
rect 26007 6502 26037 6554
rect 26037 6502 26049 6554
rect 26049 6502 26063 6554
rect 26087 6502 26101 6554
rect 26101 6502 26113 6554
rect 26113 6502 26143 6554
rect 26167 6502 26177 6554
rect 26177 6502 26223 6554
rect 25927 6500 25983 6502
rect 26007 6500 26063 6502
rect 26087 6500 26143 6502
rect 26167 6500 26223 6502
rect 28538 6196 28540 6216
rect 28540 6196 28592 6216
rect 28592 6196 28594 6216
rect 28538 6160 28594 6196
rect 25927 5466 25983 5468
rect 26007 5466 26063 5468
rect 26087 5466 26143 5468
rect 26167 5466 26223 5468
rect 25927 5414 25973 5466
rect 25973 5414 25983 5466
rect 26007 5414 26037 5466
rect 26037 5414 26049 5466
rect 26049 5414 26063 5466
rect 26087 5414 26101 5466
rect 26101 5414 26113 5466
rect 26113 5414 26143 5466
rect 26167 5414 26177 5466
rect 26177 5414 26223 5466
rect 25927 5412 25983 5414
rect 26007 5412 26063 5414
rect 26087 5412 26143 5414
rect 26167 5412 26223 5414
rect 25267 4922 25323 4924
rect 25347 4922 25403 4924
rect 25427 4922 25483 4924
rect 25507 4922 25563 4924
rect 25267 4870 25313 4922
rect 25313 4870 25323 4922
rect 25347 4870 25377 4922
rect 25377 4870 25389 4922
rect 25389 4870 25403 4922
rect 25427 4870 25441 4922
rect 25441 4870 25453 4922
rect 25453 4870 25483 4922
rect 25507 4870 25517 4922
rect 25517 4870 25563 4922
rect 25267 4868 25323 4870
rect 25347 4868 25403 4870
rect 25427 4868 25483 4870
rect 25507 4868 25563 4870
rect 25927 4378 25983 4380
rect 26007 4378 26063 4380
rect 26087 4378 26143 4380
rect 26167 4378 26223 4380
rect 25927 4326 25973 4378
rect 25973 4326 25983 4378
rect 26007 4326 26037 4378
rect 26037 4326 26049 4378
rect 26049 4326 26063 4378
rect 26087 4326 26101 4378
rect 26101 4326 26113 4378
rect 26113 4326 26143 4378
rect 26167 4326 26177 4378
rect 26177 4326 26223 4378
rect 25927 4324 25983 4326
rect 26007 4324 26063 4326
rect 26087 4324 26143 4326
rect 26167 4324 26223 4326
rect 25267 3834 25323 3836
rect 25347 3834 25403 3836
rect 25427 3834 25483 3836
rect 25507 3834 25563 3836
rect 25267 3782 25313 3834
rect 25313 3782 25323 3834
rect 25347 3782 25377 3834
rect 25377 3782 25389 3834
rect 25389 3782 25403 3834
rect 25427 3782 25441 3834
rect 25441 3782 25453 3834
rect 25453 3782 25483 3834
rect 25507 3782 25517 3834
rect 25517 3782 25563 3834
rect 25267 3780 25323 3782
rect 25347 3780 25403 3782
rect 25427 3780 25483 3782
rect 25507 3780 25563 3782
rect 25927 3290 25983 3292
rect 26007 3290 26063 3292
rect 26087 3290 26143 3292
rect 26167 3290 26223 3292
rect 25927 3238 25973 3290
rect 25973 3238 25983 3290
rect 26007 3238 26037 3290
rect 26037 3238 26049 3290
rect 26049 3238 26063 3290
rect 26087 3238 26101 3290
rect 26101 3238 26113 3290
rect 26113 3238 26143 3290
rect 26167 3238 26177 3290
rect 26177 3238 26223 3290
rect 25927 3236 25983 3238
rect 26007 3236 26063 3238
rect 26087 3236 26143 3238
rect 26167 3236 26223 3238
rect 25267 2746 25323 2748
rect 25347 2746 25403 2748
rect 25427 2746 25483 2748
rect 25507 2746 25563 2748
rect 25267 2694 25313 2746
rect 25313 2694 25323 2746
rect 25347 2694 25377 2746
rect 25377 2694 25389 2746
rect 25389 2694 25403 2746
rect 25427 2694 25441 2746
rect 25441 2694 25453 2746
rect 25453 2694 25483 2746
rect 25507 2694 25517 2746
rect 25517 2694 25563 2746
rect 25267 2692 25323 2694
rect 25347 2692 25403 2694
rect 25427 2692 25483 2694
rect 25507 2692 25563 2694
rect 18981 2202 19037 2204
rect 19061 2202 19117 2204
rect 19141 2202 19197 2204
rect 19221 2202 19277 2204
rect 18981 2150 19027 2202
rect 19027 2150 19037 2202
rect 19061 2150 19091 2202
rect 19091 2150 19103 2202
rect 19103 2150 19117 2202
rect 19141 2150 19155 2202
rect 19155 2150 19167 2202
rect 19167 2150 19197 2202
rect 19221 2150 19231 2202
rect 19231 2150 19277 2202
rect 18981 2148 19037 2150
rect 19061 2148 19117 2150
rect 19141 2148 19197 2150
rect 19221 2148 19277 2150
rect 25927 2202 25983 2204
rect 26007 2202 26063 2204
rect 26087 2202 26143 2204
rect 26167 2202 26223 2204
rect 25927 2150 25973 2202
rect 25973 2150 25983 2202
rect 26007 2150 26037 2202
rect 26037 2150 26049 2202
rect 26049 2150 26063 2202
rect 26087 2150 26101 2202
rect 26101 2150 26113 2202
rect 26113 2150 26143 2202
rect 26167 2150 26177 2202
rect 26177 2150 26223 2202
rect 25927 2148 25983 2150
rect 26007 2148 26063 2150
rect 26087 2148 26143 2150
rect 26167 2148 26223 2150
<< metal3 >>
rect 0 27978 800 28008
rect 0 27888 858 27978
rect 798 27706 858 27888
rect 4419 27776 4735 27777
rect 4419 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4735 27776
rect 4419 27711 4735 27712
rect 11365 27776 11681 27777
rect 11365 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11681 27776
rect 11365 27711 11681 27712
rect 18311 27776 18627 27777
rect 18311 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18627 27776
rect 18311 27711 18627 27712
rect 25257 27776 25573 27777
rect 25257 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25573 27776
rect 25257 27711 25573 27712
rect 1485 27706 1551 27709
rect 798 27704 1551 27706
rect 798 27648 1490 27704
rect 1546 27648 1551 27704
rect 798 27646 1551 27648
rect 1485 27643 1551 27646
rect 5079 27232 5395 27233
rect 5079 27168 5085 27232
rect 5149 27168 5165 27232
rect 5229 27168 5245 27232
rect 5309 27168 5325 27232
rect 5389 27168 5395 27232
rect 5079 27167 5395 27168
rect 12025 27232 12341 27233
rect 12025 27168 12031 27232
rect 12095 27168 12111 27232
rect 12175 27168 12191 27232
rect 12255 27168 12271 27232
rect 12335 27168 12341 27232
rect 12025 27167 12341 27168
rect 18971 27232 19287 27233
rect 18971 27168 18977 27232
rect 19041 27168 19057 27232
rect 19121 27168 19137 27232
rect 19201 27168 19217 27232
rect 19281 27168 19287 27232
rect 18971 27167 19287 27168
rect 25917 27232 26233 27233
rect 25917 27168 25923 27232
rect 25987 27168 26003 27232
rect 26067 27168 26083 27232
rect 26147 27168 26163 27232
rect 26227 27168 26233 27232
rect 25917 27167 26233 27168
rect 4419 26688 4735 26689
rect 4419 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4735 26688
rect 4419 26623 4735 26624
rect 11365 26688 11681 26689
rect 11365 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11681 26688
rect 11365 26623 11681 26624
rect 18311 26688 18627 26689
rect 18311 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18627 26688
rect 18311 26623 18627 26624
rect 25257 26688 25573 26689
rect 25257 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25573 26688
rect 25257 26623 25573 26624
rect 5079 26144 5395 26145
rect 5079 26080 5085 26144
rect 5149 26080 5165 26144
rect 5229 26080 5245 26144
rect 5309 26080 5325 26144
rect 5389 26080 5395 26144
rect 5079 26079 5395 26080
rect 12025 26144 12341 26145
rect 12025 26080 12031 26144
rect 12095 26080 12111 26144
rect 12175 26080 12191 26144
rect 12255 26080 12271 26144
rect 12335 26080 12341 26144
rect 12025 26079 12341 26080
rect 18971 26144 19287 26145
rect 18971 26080 18977 26144
rect 19041 26080 19057 26144
rect 19121 26080 19137 26144
rect 19201 26080 19217 26144
rect 19281 26080 19287 26144
rect 18971 26079 19287 26080
rect 25917 26144 26233 26145
rect 25917 26080 25923 26144
rect 25987 26080 26003 26144
rect 26067 26080 26083 26144
rect 26147 26080 26163 26144
rect 26227 26080 26233 26144
rect 25917 26079 26233 26080
rect 4419 25600 4735 25601
rect 4419 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4735 25600
rect 4419 25535 4735 25536
rect 11365 25600 11681 25601
rect 11365 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11681 25600
rect 11365 25535 11681 25536
rect 18311 25600 18627 25601
rect 18311 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18627 25600
rect 18311 25535 18627 25536
rect 25257 25600 25573 25601
rect 25257 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25573 25600
rect 25257 25535 25573 25536
rect 28533 25258 28599 25261
rect 29200 25258 30000 25288
rect 28533 25256 30000 25258
rect 28533 25200 28538 25256
rect 28594 25200 30000 25256
rect 28533 25198 30000 25200
rect 28533 25195 28599 25198
rect 29200 25168 30000 25198
rect 5079 25056 5395 25057
rect 5079 24992 5085 25056
rect 5149 24992 5165 25056
rect 5229 24992 5245 25056
rect 5309 24992 5325 25056
rect 5389 24992 5395 25056
rect 5079 24991 5395 24992
rect 12025 25056 12341 25057
rect 12025 24992 12031 25056
rect 12095 24992 12111 25056
rect 12175 24992 12191 25056
rect 12255 24992 12271 25056
rect 12335 24992 12341 25056
rect 12025 24991 12341 24992
rect 18971 25056 19287 25057
rect 18971 24992 18977 25056
rect 19041 24992 19057 25056
rect 19121 24992 19137 25056
rect 19201 24992 19217 25056
rect 19281 24992 19287 25056
rect 18971 24991 19287 24992
rect 25917 25056 26233 25057
rect 25917 24992 25923 25056
rect 25987 24992 26003 25056
rect 26067 24992 26083 25056
rect 26147 24992 26163 25056
rect 26227 24992 26233 25056
rect 25917 24991 26233 24992
rect 4419 24512 4735 24513
rect 4419 24448 4425 24512
rect 4489 24448 4505 24512
rect 4569 24448 4585 24512
rect 4649 24448 4665 24512
rect 4729 24448 4735 24512
rect 4419 24447 4735 24448
rect 11365 24512 11681 24513
rect 11365 24448 11371 24512
rect 11435 24448 11451 24512
rect 11515 24448 11531 24512
rect 11595 24448 11611 24512
rect 11675 24448 11681 24512
rect 11365 24447 11681 24448
rect 18311 24512 18627 24513
rect 18311 24448 18317 24512
rect 18381 24448 18397 24512
rect 18461 24448 18477 24512
rect 18541 24448 18557 24512
rect 18621 24448 18627 24512
rect 18311 24447 18627 24448
rect 25257 24512 25573 24513
rect 25257 24448 25263 24512
rect 25327 24448 25343 24512
rect 25407 24448 25423 24512
rect 25487 24448 25503 24512
rect 25567 24448 25573 24512
rect 25257 24447 25573 24448
rect 5079 23968 5395 23969
rect 5079 23904 5085 23968
rect 5149 23904 5165 23968
rect 5229 23904 5245 23968
rect 5309 23904 5325 23968
rect 5389 23904 5395 23968
rect 5079 23903 5395 23904
rect 12025 23968 12341 23969
rect 12025 23904 12031 23968
rect 12095 23904 12111 23968
rect 12175 23904 12191 23968
rect 12255 23904 12271 23968
rect 12335 23904 12341 23968
rect 12025 23903 12341 23904
rect 18971 23968 19287 23969
rect 18971 23904 18977 23968
rect 19041 23904 19057 23968
rect 19121 23904 19137 23968
rect 19201 23904 19217 23968
rect 19281 23904 19287 23968
rect 18971 23903 19287 23904
rect 25917 23968 26233 23969
rect 25917 23904 25923 23968
rect 25987 23904 26003 23968
rect 26067 23904 26083 23968
rect 26147 23904 26163 23968
rect 26227 23904 26233 23968
rect 25917 23903 26233 23904
rect 4419 23424 4735 23425
rect 4419 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4735 23424
rect 4419 23359 4735 23360
rect 11365 23424 11681 23425
rect 11365 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11681 23424
rect 11365 23359 11681 23360
rect 18311 23424 18627 23425
rect 18311 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18627 23424
rect 18311 23359 18627 23360
rect 25257 23424 25573 23425
rect 25257 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25573 23424
rect 25257 23359 25573 23360
rect 5079 22880 5395 22881
rect 5079 22816 5085 22880
rect 5149 22816 5165 22880
rect 5229 22816 5245 22880
rect 5309 22816 5325 22880
rect 5389 22816 5395 22880
rect 5079 22815 5395 22816
rect 12025 22880 12341 22881
rect 12025 22816 12031 22880
rect 12095 22816 12111 22880
rect 12175 22816 12191 22880
rect 12255 22816 12271 22880
rect 12335 22816 12341 22880
rect 12025 22815 12341 22816
rect 18971 22880 19287 22881
rect 18971 22816 18977 22880
rect 19041 22816 19057 22880
rect 19121 22816 19137 22880
rect 19201 22816 19217 22880
rect 19281 22816 19287 22880
rect 18971 22815 19287 22816
rect 25917 22880 26233 22881
rect 25917 22816 25923 22880
rect 25987 22816 26003 22880
rect 26067 22816 26083 22880
rect 26147 22816 26163 22880
rect 26227 22816 26233 22880
rect 25917 22815 26233 22816
rect 4419 22336 4735 22337
rect 4419 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4735 22336
rect 4419 22271 4735 22272
rect 11365 22336 11681 22337
rect 11365 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11681 22336
rect 11365 22271 11681 22272
rect 18311 22336 18627 22337
rect 18311 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18627 22336
rect 18311 22271 18627 22272
rect 25257 22336 25573 22337
rect 25257 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25573 22336
rect 25257 22271 25573 22272
rect 5079 21792 5395 21793
rect 5079 21728 5085 21792
rect 5149 21728 5165 21792
rect 5229 21728 5245 21792
rect 5309 21728 5325 21792
rect 5389 21728 5395 21792
rect 5079 21727 5395 21728
rect 12025 21792 12341 21793
rect 12025 21728 12031 21792
rect 12095 21728 12111 21792
rect 12175 21728 12191 21792
rect 12255 21728 12271 21792
rect 12335 21728 12341 21792
rect 12025 21727 12341 21728
rect 18971 21792 19287 21793
rect 18971 21728 18977 21792
rect 19041 21728 19057 21792
rect 19121 21728 19137 21792
rect 19201 21728 19217 21792
rect 19281 21728 19287 21792
rect 18971 21727 19287 21728
rect 25917 21792 26233 21793
rect 25917 21728 25923 21792
rect 25987 21728 26003 21792
rect 26067 21728 26083 21792
rect 26147 21728 26163 21792
rect 26227 21728 26233 21792
rect 25917 21727 26233 21728
rect 4419 21248 4735 21249
rect 4419 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4735 21248
rect 4419 21183 4735 21184
rect 11365 21248 11681 21249
rect 11365 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11681 21248
rect 11365 21183 11681 21184
rect 18311 21248 18627 21249
rect 18311 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18627 21248
rect 18311 21183 18627 21184
rect 25257 21248 25573 21249
rect 25257 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25573 21248
rect 25257 21183 25573 21184
rect 5079 20704 5395 20705
rect 5079 20640 5085 20704
rect 5149 20640 5165 20704
rect 5229 20640 5245 20704
rect 5309 20640 5325 20704
rect 5389 20640 5395 20704
rect 5079 20639 5395 20640
rect 12025 20704 12341 20705
rect 12025 20640 12031 20704
rect 12095 20640 12111 20704
rect 12175 20640 12191 20704
rect 12255 20640 12271 20704
rect 12335 20640 12341 20704
rect 12025 20639 12341 20640
rect 18971 20704 19287 20705
rect 18971 20640 18977 20704
rect 19041 20640 19057 20704
rect 19121 20640 19137 20704
rect 19201 20640 19217 20704
rect 19281 20640 19287 20704
rect 18971 20639 19287 20640
rect 25917 20704 26233 20705
rect 25917 20640 25923 20704
rect 25987 20640 26003 20704
rect 26067 20640 26083 20704
rect 26147 20640 26163 20704
rect 26227 20640 26233 20704
rect 25917 20639 26233 20640
rect 4419 20160 4735 20161
rect 4419 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4735 20160
rect 4419 20095 4735 20096
rect 11365 20160 11681 20161
rect 11365 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11681 20160
rect 11365 20095 11681 20096
rect 18311 20160 18627 20161
rect 18311 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18627 20160
rect 18311 20095 18627 20096
rect 25257 20160 25573 20161
rect 25257 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25573 20160
rect 25257 20095 25573 20096
rect 5079 19616 5395 19617
rect 5079 19552 5085 19616
rect 5149 19552 5165 19616
rect 5229 19552 5245 19616
rect 5309 19552 5325 19616
rect 5389 19552 5395 19616
rect 5079 19551 5395 19552
rect 12025 19616 12341 19617
rect 12025 19552 12031 19616
rect 12095 19552 12111 19616
rect 12175 19552 12191 19616
rect 12255 19552 12271 19616
rect 12335 19552 12341 19616
rect 12025 19551 12341 19552
rect 18971 19616 19287 19617
rect 18971 19552 18977 19616
rect 19041 19552 19057 19616
rect 19121 19552 19137 19616
rect 19201 19552 19217 19616
rect 19281 19552 19287 19616
rect 18971 19551 19287 19552
rect 25917 19616 26233 19617
rect 25917 19552 25923 19616
rect 25987 19552 26003 19616
rect 26067 19552 26083 19616
rect 26147 19552 26163 19616
rect 26227 19552 26233 19616
rect 25917 19551 26233 19552
rect 4419 19072 4735 19073
rect 4419 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4735 19072
rect 4419 19007 4735 19008
rect 11365 19072 11681 19073
rect 11365 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11681 19072
rect 11365 19007 11681 19008
rect 18311 19072 18627 19073
rect 18311 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18627 19072
rect 18311 19007 18627 19008
rect 25257 19072 25573 19073
rect 25257 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25573 19072
rect 25257 19007 25573 19008
rect 5079 18528 5395 18529
rect 0 18458 800 18488
rect 5079 18464 5085 18528
rect 5149 18464 5165 18528
rect 5229 18464 5245 18528
rect 5309 18464 5325 18528
rect 5389 18464 5395 18528
rect 5079 18463 5395 18464
rect 12025 18528 12341 18529
rect 12025 18464 12031 18528
rect 12095 18464 12111 18528
rect 12175 18464 12191 18528
rect 12255 18464 12271 18528
rect 12335 18464 12341 18528
rect 12025 18463 12341 18464
rect 18971 18528 19287 18529
rect 18971 18464 18977 18528
rect 19041 18464 19057 18528
rect 19121 18464 19137 18528
rect 19201 18464 19217 18528
rect 19281 18464 19287 18528
rect 18971 18463 19287 18464
rect 25917 18528 26233 18529
rect 25917 18464 25923 18528
rect 25987 18464 26003 18528
rect 26067 18464 26083 18528
rect 26147 18464 26163 18528
rect 26227 18464 26233 18528
rect 25917 18463 26233 18464
rect 933 18458 999 18461
rect 0 18456 999 18458
rect 0 18400 938 18456
rect 994 18400 999 18456
rect 0 18398 999 18400
rect 0 18368 800 18398
rect 933 18395 999 18398
rect 4419 17984 4735 17985
rect 4419 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4735 17984
rect 4419 17919 4735 17920
rect 11365 17984 11681 17985
rect 11365 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11681 17984
rect 11365 17919 11681 17920
rect 18311 17984 18627 17985
rect 18311 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18627 17984
rect 18311 17919 18627 17920
rect 25257 17984 25573 17985
rect 25257 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25573 17984
rect 25257 17919 25573 17920
rect 5079 17440 5395 17441
rect 5079 17376 5085 17440
rect 5149 17376 5165 17440
rect 5229 17376 5245 17440
rect 5309 17376 5325 17440
rect 5389 17376 5395 17440
rect 5079 17375 5395 17376
rect 12025 17440 12341 17441
rect 12025 17376 12031 17440
rect 12095 17376 12111 17440
rect 12175 17376 12191 17440
rect 12255 17376 12271 17440
rect 12335 17376 12341 17440
rect 12025 17375 12341 17376
rect 18971 17440 19287 17441
rect 18971 17376 18977 17440
rect 19041 17376 19057 17440
rect 19121 17376 19137 17440
rect 19201 17376 19217 17440
rect 19281 17376 19287 17440
rect 18971 17375 19287 17376
rect 25917 17440 26233 17441
rect 25917 17376 25923 17440
rect 25987 17376 26003 17440
rect 26067 17376 26083 17440
rect 26147 17376 26163 17440
rect 26227 17376 26233 17440
rect 25917 17375 26233 17376
rect 4419 16896 4735 16897
rect 4419 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4735 16896
rect 4419 16831 4735 16832
rect 11365 16896 11681 16897
rect 11365 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11681 16896
rect 11365 16831 11681 16832
rect 18311 16896 18627 16897
rect 18311 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18627 16896
rect 18311 16831 18627 16832
rect 25257 16896 25573 16897
rect 25257 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25573 16896
rect 25257 16831 25573 16832
rect 5079 16352 5395 16353
rect 5079 16288 5085 16352
rect 5149 16288 5165 16352
rect 5229 16288 5245 16352
rect 5309 16288 5325 16352
rect 5389 16288 5395 16352
rect 5079 16287 5395 16288
rect 12025 16352 12341 16353
rect 12025 16288 12031 16352
rect 12095 16288 12111 16352
rect 12175 16288 12191 16352
rect 12255 16288 12271 16352
rect 12335 16288 12341 16352
rect 12025 16287 12341 16288
rect 18971 16352 19287 16353
rect 18971 16288 18977 16352
rect 19041 16288 19057 16352
rect 19121 16288 19137 16352
rect 19201 16288 19217 16352
rect 19281 16288 19287 16352
rect 18971 16287 19287 16288
rect 25917 16352 26233 16353
rect 25917 16288 25923 16352
rect 25987 16288 26003 16352
rect 26067 16288 26083 16352
rect 26147 16288 26163 16352
rect 26227 16288 26233 16352
rect 25917 16287 26233 16288
rect 4419 15808 4735 15809
rect 4419 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4735 15808
rect 4419 15743 4735 15744
rect 11365 15808 11681 15809
rect 11365 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11681 15808
rect 11365 15743 11681 15744
rect 18311 15808 18627 15809
rect 18311 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18627 15808
rect 18311 15743 18627 15744
rect 25257 15808 25573 15809
rect 25257 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25573 15808
rect 25257 15743 25573 15744
rect 24894 15676 24900 15740
rect 24964 15676 24970 15740
rect 29200 15738 30000 15768
rect 26190 15678 30000 15738
rect 24902 15602 24962 15676
rect 26190 15602 26250 15678
rect 29200 15648 30000 15678
rect 24902 15542 26250 15602
rect 5079 15264 5395 15265
rect 5079 15200 5085 15264
rect 5149 15200 5165 15264
rect 5229 15200 5245 15264
rect 5309 15200 5325 15264
rect 5389 15200 5395 15264
rect 5079 15199 5395 15200
rect 12025 15264 12341 15265
rect 12025 15200 12031 15264
rect 12095 15200 12111 15264
rect 12175 15200 12191 15264
rect 12255 15200 12271 15264
rect 12335 15200 12341 15264
rect 12025 15199 12341 15200
rect 18971 15264 19287 15265
rect 18971 15200 18977 15264
rect 19041 15200 19057 15264
rect 19121 15200 19137 15264
rect 19201 15200 19217 15264
rect 19281 15200 19287 15264
rect 18971 15199 19287 15200
rect 25917 15264 26233 15265
rect 25917 15200 25923 15264
rect 25987 15200 26003 15264
rect 26067 15200 26083 15264
rect 26147 15200 26163 15264
rect 26227 15200 26233 15264
rect 25917 15199 26233 15200
rect 4419 14720 4735 14721
rect 4419 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4735 14720
rect 4419 14655 4735 14656
rect 11365 14720 11681 14721
rect 11365 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11681 14720
rect 11365 14655 11681 14656
rect 18311 14720 18627 14721
rect 18311 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18627 14720
rect 18311 14655 18627 14656
rect 25257 14720 25573 14721
rect 25257 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25573 14720
rect 25257 14655 25573 14656
rect 5079 14176 5395 14177
rect 5079 14112 5085 14176
rect 5149 14112 5165 14176
rect 5229 14112 5245 14176
rect 5309 14112 5325 14176
rect 5389 14112 5395 14176
rect 5079 14111 5395 14112
rect 12025 14176 12341 14177
rect 12025 14112 12031 14176
rect 12095 14112 12111 14176
rect 12175 14112 12191 14176
rect 12255 14112 12271 14176
rect 12335 14112 12341 14176
rect 12025 14111 12341 14112
rect 18971 14176 19287 14177
rect 18971 14112 18977 14176
rect 19041 14112 19057 14176
rect 19121 14112 19137 14176
rect 19201 14112 19217 14176
rect 19281 14112 19287 14176
rect 18971 14111 19287 14112
rect 25917 14176 26233 14177
rect 25917 14112 25923 14176
rect 25987 14112 26003 14176
rect 26067 14112 26083 14176
rect 26147 14112 26163 14176
rect 26227 14112 26233 14176
rect 25917 14111 26233 14112
rect 4419 13632 4735 13633
rect 4419 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4735 13632
rect 4419 13567 4735 13568
rect 11365 13632 11681 13633
rect 11365 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11681 13632
rect 11365 13567 11681 13568
rect 18311 13632 18627 13633
rect 18311 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18627 13632
rect 18311 13567 18627 13568
rect 25257 13632 25573 13633
rect 25257 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25573 13632
rect 25257 13567 25573 13568
rect 5079 13088 5395 13089
rect 5079 13024 5085 13088
rect 5149 13024 5165 13088
rect 5229 13024 5245 13088
rect 5309 13024 5325 13088
rect 5389 13024 5395 13088
rect 5079 13023 5395 13024
rect 12025 13088 12341 13089
rect 12025 13024 12031 13088
rect 12095 13024 12111 13088
rect 12175 13024 12191 13088
rect 12255 13024 12271 13088
rect 12335 13024 12341 13088
rect 12025 13023 12341 13024
rect 18971 13088 19287 13089
rect 18971 13024 18977 13088
rect 19041 13024 19057 13088
rect 19121 13024 19137 13088
rect 19201 13024 19217 13088
rect 19281 13024 19287 13088
rect 18971 13023 19287 13024
rect 25917 13088 26233 13089
rect 25917 13024 25923 13088
rect 25987 13024 26003 13088
rect 26067 13024 26083 13088
rect 26147 13024 26163 13088
rect 26227 13024 26233 13088
rect 25917 13023 26233 13024
rect 4419 12544 4735 12545
rect 4419 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4735 12544
rect 4419 12479 4735 12480
rect 11365 12544 11681 12545
rect 11365 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11681 12544
rect 11365 12479 11681 12480
rect 18311 12544 18627 12545
rect 18311 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18627 12544
rect 18311 12479 18627 12480
rect 25257 12544 25573 12545
rect 25257 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25573 12544
rect 25257 12479 25573 12480
rect 5079 12000 5395 12001
rect 5079 11936 5085 12000
rect 5149 11936 5165 12000
rect 5229 11936 5245 12000
rect 5309 11936 5325 12000
rect 5389 11936 5395 12000
rect 5079 11935 5395 11936
rect 12025 12000 12341 12001
rect 12025 11936 12031 12000
rect 12095 11936 12111 12000
rect 12175 11936 12191 12000
rect 12255 11936 12271 12000
rect 12335 11936 12341 12000
rect 12025 11935 12341 11936
rect 18971 12000 19287 12001
rect 18971 11936 18977 12000
rect 19041 11936 19057 12000
rect 19121 11936 19137 12000
rect 19201 11936 19217 12000
rect 19281 11936 19287 12000
rect 18971 11935 19287 11936
rect 25917 12000 26233 12001
rect 25917 11936 25923 12000
rect 25987 11936 26003 12000
rect 26067 11936 26083 12000
rect 26147 11936 26163 12000
rect 26227 11936 26233 12000
rect 25917 11935 26233 11936
rect 4419 11456 4735 11457
rect 4419 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4735 11456
rect 4419 11391 4735 11392
rect 11365 11456 11681 11457
rect 11365 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11681 11456
rect 11365 11391 11681 11392
rect 18311 11456 18627 11457
rect 18311 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18627 11456
rect 18311 11391 18627 11392
rect 25257 11456 25573 11457
rect 25257 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25573 11456
rect 25257 11391 25573 11392
rect 5079 10912 5395 10913
rect 5079 10848 5085 10912
rect 5149 10848 5165 10912
rect 5229 10848 5245 10912
rect 5309 10848 5325 10912
rect 5389 10848 5395 10912
rect 5079 10847 5395 10848
rect 12025 10912 12341 10913
rect 12025 10848 12031 10912
rect 12095 10848 12111 10912
rect 12175 10848 12191 10912
rect 12255 10848 12271 10912
rect 12335 10848 12341 10912
rect 12025 10847 12341 10848
rect 18971 10912 19287 10913
rect 18971 10848 18977 10912
rect 19041 10848 19057 10912
rect 19121 10848 19137 10912
rect 19201 10848 19217 10912
rect 19281 10848 19287 10912
rect 18971 10847 19287 10848
rect 25917 10912 26233 10913
rect 25917 10848 25923 10912
rect 25987 10848 26003 10912
rect 26067 10848 26083 10912
rect 26147 10848 26163 10912
rect 26227 10848 26233 10912
rect 25917 10847 26233 10848
rect 4419 10368 4735 10369
rect 4419 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4735 10368
rect 4419 10303 4735 10304
rect 11365 10368 11681 10369
rect 11365 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11681 10368
rect 11365 10303 11681 10304
rect 18311 10368 18627 10369
rect 18311 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18627 10368
rect 18311 10303 18627 10304
rect 25257 10368 25573 10369
rect 25257 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25573 10368
rect 25257 10303 25573 10304
rect 5079 9824 5395 9825
rect 5079 9760 5085 9824
rect 5149 9760 5165 9824
rect 5229 9760 5245 9824
rect 5309 9760 5325 9824
rect 5389 9760 5395 9824
rect 5079 9759 5395 9760
rect 12025 9824 12341 9825
rect 12025 9760 12031 9824
rect 12095 9760 12111 9824
rect 12175 9760 12191 9824
rect 12255 9760 12271 9824
rect 12335 9760 12341 9824
rect 12025 9759 12341 9760
rect 18971 9824 19287 9825
rect 18971 9760 18977 9824
rect 19041 9760 19057 9824
rect 19121 9760 19137 9824
rect 19201 9760 19217 9824
rect 19281 9760 19287 9824
rect 18971 9759 19287 9760
rect 25917 9824 26233 9825
rect 25917 9760 25923 9824
rect 25987 9760 26003 9824
rect 26067 9760 26083 9824
rect 26147 9760 26163 9824
rect 26227 9760 26233 9824
rect 25917 9759 26233 9760
rect 17769 9482 17835 9485
rect 17726 9480 17835 9482
rect 17726 9424 17774 9480
rect 17830 9424 17835 9480
rect 17726 9419 17835 9424
rect 17726 9349 17786 9419
rect 17726 9344 17835 9349
rect 17726 9288 17774 9344
rect 17830 9288 17835 9344
rect 17726 9286 17835 9288
rect 17769 9283 17835 9286
rect 4419 9280 4735 9281
rect 4419 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4735 9280
rect 4419 9215 4735 9216
rect 11365 9280 11681 9281
rect 11365 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11681 9280
rect 11365 9215 11681 9216
rect 18311 9280 18627 9281
rect 18311 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18627 9280
rect 18311 9215 18627 9216
rect 25257 9280 25573 9281
rect 25257 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25573 9280
rect 25257 9215 25573 9216
rect 16757 9074 16823 9077
rect 18873 9074 18939 9077
rect 16757 9072 18939 9074
rect 16757 9016 16762 9072
rect 16818 9016 18878 9072
rect 18934 9016 18939 9072
rect 16757 9014 18939 9016
rect 16757 9011 16823 9014
rect 18873 9011 18939 9014
rect 0 8938 800 8968
rect 933 8938 999 8941
rect 0 8936 999 8938
rect 0 8880 938 8936
rect 994 8880 999 8936
rect 0 8878 999 8880
rect 0 8848 800 8878
rect 933 8875 999 8878
rect 5079 8736 5395 8737
rect 5079 8672 5085 8736
rect 5149 8672 5165 8736
rect 5229 8672 5245 8736
rect 5309 8672 5325 8736
rect 5389 8672 5395 8736
rect 5079 8671 5395 8672
rect 12025 8736 12341 8737
rect 12025 8672 12031 8736
rect 12095 8672 12111 8736
rect 12175 8672 12191 8736
rect 12255 8672 12271 8736
rect 12335 8672 12341 8736
rect 12025 8671 12341 8672
rect 18971 8736 19287 8737
rect 18971 8672 18977 8736
rect 19041 8672 19057 8736
rect 19121 8672 19137 8736
rect 19201 8672 19217 8736
rect 19281 8672 19287 8736
rect 18971 8671 19287 8672
rect 25917 8736 26233 8737
rect 25917 8672 25923 8736
rect 25987 8672 26003 8736
rect 26067 8672 26083 8736
rect 26147 8672 26163 8736
rect 26227 8672 26233 8736
rect 25917 8671 26233 8672
rect 21817 8258 21883 8261
rect 24894 8258 24900 8260
rect 21817 8256 24900 8258
rect 21817 8200 21822 8256
rect 21878 8200 24900 8256
rect 21817 8198 24900 8200
rect 21817 8195 21883 8198
rect 24894 8196 24900 8198
rect 24964 8196 24970 8260
rect 4419 8192 4735 8193
rect 4419 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4735 8192
rect 4419 8127 4735 8128
rect 11365 8192 11681 8193
rect 11365 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11681 8192
rect 11365 8127 11681 8128
rect 18311 8192 18627 8193
rect 18311 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18627 8192
rect 18311 8127 18627 8128
rect 25257 8192 25573 8193
rect 25257 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25573 8192
rect 25257 8127 25573 8128
rect 17769 7850 17835 7853
rect 18689 7850 18755 7853
rect 17769 7848 18755 7850
rect 17769 7792 17774 7848
rect 17830 7792 18694 7848
rect 18750 7792 18755 7848
rect 17769 7790 18755 7792
rect 17769 7787 17835 7790
rect 18689 7787 18755 7790
rect 5079 7648 5395 7649
rect 5079 7584 5085 7648
rect 5149 7584 5165 7648
rect 5229 7584 5245 7648
rect 5309 7584 5325 7648
rect 5389 7584 5395 7648
rect 5079 7583 5395 7584
rect 12025 7648 12341 7649
rect 12025 7584 12031 7648
rect 12095 7584 12111 7648
rect 12175 7584 12191 7648
rect 12255 7584 12271 7648
rect 12335 7584 12341 7648
rect 12025 7583 12341 7584
rect 18971 7648 19287 7649
rect 18971 7584 18977 7648
rect 19041 7584 19057 7648
rect 19121 7584 19137 7648
rect 19201 7584 19217 7648
rect 19281 7584 19287 7648
rect 18971 7583 19287 7584
rect 25917 7648 26233 7649
rect 25917 7584 25923 7648
rect 25987 7584 26003 7648
rect 26067 7584 26083 7648
rect 26147 7584 26163 7648
rect 26227 7584 26233 7648
rect 25917 7583 26233 7584
rect 17861 7306 17927 7309
rect 20805 7306 20871 7309
rect 17861 7304 20871 7306
rect 17861 7248 17866 7304
rect 17922 7248 20810 7304
rect 20866 7248 20871 7304
rect 17861 7246 20871 7248
rect 17861 7243 17927 7246
rect 20805 7243 20871 7246
rect 21909 7306 21975 7309
rect 22921 7306 22987 7309
rect 21909 7304 22987 7306
rect 21909 7248 21914 7304
rect 21970 7248 22926 7304
rect 22982 7248 22987 7304
rect 21909 7246 22987 7248
rect 21909 7243 21975 7246
rect 22921 7243 22987 7246
rect 4419 7104 4735 7105
rect 4419 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4735 7104
rect 4419 7039 4735 7040
rect 11365 7104 11681 7105
rect 11365 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11681 7104
rect 11365 7039 11681 7040
rect 18311 7104 18627 7105
rect 18311 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18627 7104
rect 18311 7039 18627 7040
rect 25257 7104 25573 7105
rect 25257 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25573 7104
rect 25257 7039 25573 7040
rect 5079 6560 5395 6561
rect 5079 6496 5085 6560
rect 5149 6496 5165 6560
rect 5229 6496 5245 6560
rect 5309 6496 5325 6560
rect 5389 6496 5395 6560
rect 5079 6495 5395 6496
rect 12025 6560 12341 6561
rect 12025 6496 12031 6560
rect 12095 6496 12111 6560
rect 12175 6496 12191 6560
rect 12255 6496 12271 6560
rect 12335 6496 12341 6560
rect 12025 6495 12341 6496
rect 18971 6560 19287 6561
rect 18971 6496 18977 6560
rect 19041 6496 19057 6560
rect 19121 6496 19137 6560
rect 19201 6496 19217 6560
rect 19281 6496 19287 6560
rect 18971 6495 19287 6496
rect 25917 6560 26233 6561
rect 25917 6496 25923 6560
rect 25987 6496 26003 6560
rect 26067 6496 26083 6560
rect 26147 6496 26163 6560
rect 26227 6496 26233 6560
rect 25917 6495 26233 6496
rect 28533 6218 28599 6221
rect 29200 6218 30000 6248
rect 28533 6216 30000 6218
rect 28533 6160 28538 6216
rect 28594 6160 30000 6216
rect 28533 6158 30000 6160
rect 28533 6155 28599 6158
rect 29200 6128 30000 6158
rect 4419 6016 4735 6017
rect 4419 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4735 6016
rect 4419 5951 4735 5952
rect 11365 6016 11681 6017
rect 11365 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11681 6016
rect 11365 5951 11681 5952
rect 18311 6016 18627 6017
rect 18311 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18627 6016
rect 18311 5951 18627 5952
rect 25257 6016 25573 6017
rect 25257 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25573 6016
rect 25257 5951 25573 5952
rect 5079 5472 5395 5473
rect 5079 5408 5085 5472
rect 5149 5408 5165 5472
rect 5229 5408 5245 5472
rect 5309 5408 5325 5472
rect 5389 5408 5395 5472
rect 5079 5407 5395 5408
rect 12025 5472 12341 5473
rect 12025 5408 12031 5472
rect 12095 5408 12111 5472
rect 12175 5408 12191 5472
rect 12255 5408 12271 5472
rect 12335 5408 12341 5472
rect 12025 5407 12341 5408
rect 18971 5472 19287 5473
rect 18971 5408 18977 5472
rect 19041 5408 19057 5472
rect 19121 5408 19137 5472
rect 19201 5408 19217 5472
rect 19281 5408 19287 5472
rect 18971 5407 19287 5408
rect 25917 5472 26233 5473
rect 25917 5408 25923 5472
rect 25987 5408 26003 5472
rect 26067 5408 26083 5472
rect 26147 5408 26163 5472
rect 26227 5408 26233 5472
rect 25917 5407 26233 5408
rect 4419 4928 4735 4929
rect 4419 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4735 4928
rect 4419 4863 4735 4864
rect 11365 4928 11681 4929
rect 11365 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11681 4928
rect 11365 4863 11681 4864
rect 18311 4928 18627 4929
rect 18311 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18627 4928
rect 18311 4863 18627 4864
rect 25257 4928 25573 4929
rect 25257 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25573 4928
rect 25257 4863 25573 4864
rect 5079 4384 5395 4385
rect 5079 4320 5085 4384
rect 5149 4320 5165 4384
rect 5229 4320 5245 4384
rect 5309 4320 5325 4384
rect 5389 4320 5395 4384
rect 5079 4319 5395 4320
rect 12025 4384 12341 4385
rect 12025 4320 12031 4384
rect 12095 4320 12111 4384
rect 12175 4320 12191 4384
rect 12255 4320 12271 4384
rect 12335 4320 12341 4384
rect 12025 4319 12341 4320
rect 18971 4384 19287 4385
rect 18971 4320 18977 4384
rect 19041 4320 19057 4384
rect 19121 4320 19137 4384
rect 19201 4320 19217 4384
rect 19281 4320 19287 4384
rect 18971 4319 19287 4320
rect 25917 4384 26233 4385
rect 25917 4320 25923 4384
rect 25987 4320 26003 4384
rect 26067 4320 26083 4384
rect 26147 4320 26163 4384
rect 26227 4320 26233 4384
rect 25917 4319 26233 4320
rect 17125 4178 17191 4181
rect 18965 4178 19031 4181
rect 17125 4176 19031 4178
rect 17125 4120 17130 4176
rect 17186 4120 18970 4176
rect 19026 4120 19031 4176
rect 17125 4118 19031 4120
rect 17125 4115 17191 4118
rect 18965 4115 19031 4118
rect 4419 3840 4735 3841
rect 4419 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4735 3840
rect 4419 3775 4735 3776
rect 11365 3840 11681 3841
rect 11365 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11681 3840
rect 11365 3775 11681 3776
rect 18311 3840 18627 3841
rect 18311 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18627 3840
rect 18311 3775 18627 3776
rect 25257 3840 25573 3841
rect 25257 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25573 3840
rect 25257 3775 25573 3776
rect 5079 3296 5395 3297
rect 5079 3232 5085 3296
rect 5149 3232 5165 3296
rect 5229 3232 5245 3296
rect 5309 3232 5325 3296
rect 5389 3232 5395 3296
rect 5079 3231 5395 3232
rect 12025 3296 12341 3297
rect 12025 3232 12031 3296
rect 12095 3232 12111 3296
rect 12175 3232 12191 3296
rect 12255 3232 12271 3296
rect 12335 3232 12341 3296
rect 12025 3231 12341 3232
rect 18971 3296 19287 3297
rect 18971 3232 18977 3296
rect 19041 3232 19057 3296
rect 19121 3232 19137 3296
rect 19201 3232 19217 3296
rect 19281 3232 19287 3296
rect 18971 3231 19287 3232
rect 25917 3296 26233 3297
rect 25917 3232 25923 3296
rect 25987 3232 26003 3296
rect 26067 3232 26083 3296
rect 26147 3232 26163 3296
rect 26227 3232 26233 3296
rect 25917 3231 26233 3232
rect 4419 2752 4735 2753
rect 4419 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4735 2752
rect 4419 2687 4735 2688
rect 11365 2752 11681 2753
rect 11365 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11681 2752
rect 11365 2687 11681 2688
rect 18311 2752 18627 2753
rect 18311 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18627 2752
rect 18311 2687 18627 2688
rect 25257 2752 25573 2753
rect 25257 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25573 2752
rect 25257 2687 25573 2688
rect 5079 2208 5395 2209
rect 5079 2144 5085 2208
rect 5149 2144 5165 2208
rect 5229 2144 5245 2208
rect 5309 2144 5325 2208
rect 5389 2144 5395 2208
rect 5079 2143 5395 2144
rect 12025 2208 12341 2209
rect 12025 2144 12031 2208
rect 12095 2144 12111 2208
rect 12175 2144 12191 2208
rect 12255 2144 12271 2208
rect 12335 2144 12341 2208
rect 12025 2143 12341 2144
rect 18971 2208 19287 2209
rect 18971 2144 18977 2208
rect 19041 2144 19057 2208
rect 19121 2144 19137 2208
rect 19201 2144 19217 2208
rect 19281 2144 19287 2208
rect 18971 2143 19287 2144
rect 25917 2208 26233 2209
rect 25917 2144 25923 2208
rect 25987 2144 26003 2208
rect 26067 2144 26083 2208
rect 26147 2144 26163 2208
rect 26227 2144 26233 2208
rect 25917 2143 26233 2144
<< via3 >>
rect 4425 27772 4489 27776
rect 4425 27716 4429 27772
rect 4429 27716 4485 27772
rect 4485 27716 4489 27772
rect 4425 27712 4489 27716
rect 4505 27772 4569 27776
rect 4505 27716 4509 27772
rect 4509 27716 4565 27772
rect 4565 27716 4569 27772
rect 4505 27712 4569 27716
rect 4585 27772 4649 27776
rect 4585 27716 4589 27772
rect 4589 27716 4645 27772
rect 4645 27716 4649 27772
rect 4585 27712 4649 27716
rect 4665 27772 4729 27776
rect 4665 27716 4669 27772
rect 4669 27716 4725 27772
rect 4725 27716 4729 27772
rect 4665 27712 4729 27716
rect 11371 27772 11435 27776
rect 11371 27716 11375 27772
rect 11375 27716 11431 27772
rect 11431 27716 11435 27772
rect 11371 27712 11435 27716
rect 11451 27772 11515 27776
rect 11451 27716 11455 27772
rect 11455 27716 11511 27772
rect 11511 27716 11515 27772
rect 11451 27712 11515 27716
rect 11531 27772 11595 27776
rect 11531 27716 11535 27772
rect 11535 27716 11591 27772
rect 11591 27716 11595 27772
rect 11531 27712 11595 27716
rect 11611 27772 11675 27776
rect 11611 27716 11615 27772
rect 11615 27716 11671 27772
rect 11671 27716 11675 27772
rect 11611 27712 11675 27716
rect 18317 27772 18381 27776
rect 18317 27716 18321 27772
rect 18321 27716 18377 27772
rect 18377 27716 18381 27772
rect 18317 27712 18381 27716
rect 18397 27772 18461 27776
rect 18397 27716 18401 27772
rect 18401 27716 18457 27772
rect 18457 27716 18461 27772
rect 18397 27712 18461 27716
rect 18477 27772 18541 27776
rect 18477 27716 18481 27772
rect 18481 27716 18537 27772
rect 18537 27716 18541 27772
rect 18477 27712 18541 27716
rect 18557 27772 18621 27776
rect 18557 27716 18561 27772
rect 18561 27716 18617 27772
rect 18617 27716 18621 27772
rect 18557 27712 18621 27716
rect 25263 27772 25327 27776
rect 25263 27716 25267 27772
rect 25267 27716 25323 27772
rect 25323 27716 25327 27772
rect 25263 27712 25327 27716
rect 25343 27772 25407 27776
rect 25343 27716 25347 27772
rect 25347 27716 25403 27772
rect 25403 27716 25407 27772
rect 25343 27712 25407 27716
rect 25423 27772 25487 27776
rect 25423 27716 25427 27772
rect 25427 27716 25483 27772
rect 25483 27716 25487 27772
rect 25423 27712 25487 27716
rect 25503 27772 25567 27776
rect 25503 27716 25507 27772
rect 25507 27716 25563 27772
rect 25563 27716 25567 27772
rect 25503 27712 25567 27716
rect 5085 27228 5149 27232
rect 5085 27172 5089 27228
rect 5089 27172 5145 27228
rect 5145 27172 5149 27228
rect 5085 27168 5149 27172
rect 5165 27228 5229 27232
rect 5165 27172 5169 27228
rect 5169 27172 5225 27228
rect 5225 27172 5229 27228
rect 5165 27168 5229 27172
rect 5245 27228 5309 27232
rect 5245 27172 5249 27228
rect 5249 27172 5305 27228
rect 5305 27172 5309 27228
rect 5245 27168 5309 27172
rect 5325 27228 5389 27232
rect 5325 27172 5329 27228
rect 5329 27172 5385 27228
rect 5385 27172 5389 27228
rect 5325 27168 5389 27172
rect 12031 27228 12095 27232
rect 12031 27172 12035 27228
rect 12035 27172 12091 27228
rect 12091 27172 12095 27228
rect 12031 27168 12095 27172
rect 12111 27228 12175 27232
rect 12111 27172 12115 27228
rect 12115 27172 12171 27228
rect 12171 27172 12175 27228
rect 12111 27168 12175 27172
rect 12191 27228 12255 27232
rect 12191 27172 12195 27228
rect 12195 27172 12251 27228
rect 12251 27172 12255 27228
rect 12191 27168 12255 27172
rect 12271 27228 12335 27232
rect 12271 27172 12275 27228
rect 12275 27172 12331 27228
rect 12331 27172 12335 27228
rect 12271 27168 12335 27172
rect 18977 27228 19041 27232
rect 18977 27172 18981 27228
rect 18981 27172 19037 27228
rect 19037 27172 19041 27228
rect 18977 27168 19041 27172
rect 19057 27228 19121 27232
rect 19057 27172 19061 27228
rect 19061 27172 19117 27228
rect 19117 27172 19121 27228
rect 19057 27168 19121 27172
rect 19137 27228 19201 27232
rect 19137 27172 19141 27228
rect 19141 27172 19197 27228
rect 19197 27172 19201 27228
rect 19137 27168 19201 27172
rect 19217 27228 19281 27232
rect 19217 27172 19221 27228
rect 19221 27172 19277 27228
rect 19277 27172 19281 27228
rect 19217 27168 19281 27172
rect 25923 27228 25987 27232
rect 25923 27172 25927 27228
rect 25927 27172 25983 27228
rect 25983 27172 25987 27228
rect 25923 27168 25987 27172
rect 26003 27228 26067 27232
rect 26003 27172 26007 27228
rect 26007 27172 26063 27228
rect 26063 27172 26067 27228
rect 26003 27168 26067 27172
rect 26083 27228 26147 27232
rect 26083 27172 26087 27228
rect 26087 27172 26143 27228
rect 26143 27172 26147 27228
rect 26083 27168 26147 27172
rect 26163 27228 26227 27232
rect 26163 27172 26167 27228
rect 26167 27172 26223 27228
rect 26223 27172 26227 27228
rect 26163 27168 26227 27172
rect 4425 26684 4489 26688
rect 4425 26628 4429 26684
rect 4429 26628 4485 26684
rect 4485 26628 4489 26684
rect 4425 26624 4489 26628
rect 4505 26684 4569 26688
rect 4505 26628 4509 26684
rect 4509 26628 4565 26684
rect 4565 26628 4569 26684
rect 4505 26624 4569 26628
rect 4585 26684 4649 26688
rect 4585 26628 4589 26684
rect 4589 26628 4645 26684
rect 4645 26628 4649 26684
rect 4585 26624 4649 26628
rect 4665 26684 4729 26688
rect 4665 26628 4669 26684
rect 4669 26628 4725 26684
rect 4725 26628 4729 26684
rect 4665 26624 4729 26628
rect 11371 26684 11435 26688
rect 11371 26628 11375 26684
rect 11375 26628 11431 26684
rect 11431 26628 11435 26684
rect 11371 26624 11435 26628
rect 11451 26684 11515 26688
rect 11451 26628 11455 26684
rect 11455 26628 11511 26684
rect 11511 26628 11515 26684
rect 11451 26624 11515 26628
rect 11531 26684 11595 26688
rect 11531 26628 11535 26684
rect 11535 26628 11591 26684
rect 11591 26628 11595 26684
rect 11531 26624 11595 26628
rect 11611 26684 11675 26688
rect 11611 26628 11615 26684
rect 11615 26628 11671 26684
rect 11671 26628 11675 26684
rect 11611 26624 11675 26628
rect 18317 26684 18381 26688
rect 18317 26628 18321 26684
rect 18321 26628 18377 26684
rect 18377 26628 18381 26684
rect 18317 26624 18381 26628
rect 18397 26684 18461 26688
rect 18397 26628 18401 26684
rect 18401 26628 18457 26684
rect 18457 26628 18461 26684
rect 18397 26624 18461 26628
rect 18477 26684 18541 26688
rect 18477 26628 18481 26684
rect 18481 26628 18537 26684
rect 18537 26628 18541 26684
rect 18477 26624 18541 26628
rect 18557 26684 18621 26688
rect 18557 26628 18561 26684
rect 18561 26628 18617 26684
rect 18617 26628 18621 26684
rect 18557 26624 18621 26628
rect 25263 26684 25327 26688
rect 25263 26628 25267 26684
rect 25267 26628 25323 26684
rect 25323 26628 25327 26684
rect 25263 26624 25327 26628
rect 25343 26684 25407 26688
rect 25343 26628 25347 26684
rect 25347 26628 25403 26684
rect 25403 26628 25407 26684
rect 25343 26624 25407 26628
rect 25423 26684 25487 26688
rect 25423 26628 25427 26684
rect 25427 26628 25483 26684
rect 25483 26628 25487 26684
rect 25423 26624 25487 26628
rect 25503 26684 25567 26688
rect 25503 26628 25507 26684
rect 25507 26628 25563 26684
rect 25563 26628 25567 26684
rect 25503 26624 25567 26628
rect 5085 26140 5149 26144
rect 5085 26084 5089 26140
rect 5089 26084 5145 26140
rect 5145 26084 5149 26140
rect 5085 26080 5149 26084
rect 5165 26140 5229 26144
rect 5165 26084 5169 26140
rect 5169 26084 5225 26140
rect 5225 26084 5229 26140
rect 5165 26080 5229 26084
rect 5245 26140 5309 26144
rect 5245 26084 5249 26140
rect 5249 26084 5305 26140
rect 5305 26084 5309 26140
rect 5245 26080 5309 26084
rect 5325 26140 5389 26144
rect 5325 26084 5329 26140
rect 5329 26084 5385 26140
rect 5385 26084 5389 26140
rect 5325 26080 5389 26084
rect 12031 26140 12095 26144
rect 12031 26084 12035 26140
rect 12035 26084 12091 26140
rect 12091 26084 12095 26140
rect 12031 26080 12095 26084
rect 12111 26140 12175 26144
rect 12111 26084 12115 26140
rect 12115 26084 12171 26140
rect 12171 26084 12175 26140
rect 12111 26080 12175 26084
rect 12191 26140 12255 26144
rect 12191 26084 12195 26140
rect 12195 26084 12251 26140
rect 12251 26084 12255 26140
rect 12191 26080 12255 26084
rect 12271 26140 12335 26144
rect 12271 26084 12275 26140
rect 12275 26084 12331 26140
rect 12331 26084 12335 26140
rect 12271 26080 12335 26084
rect 18977 26140 19041 26144
rect 18977 26084 18981 26140
rect 18981 26084 19037 26140
rect 19037 26084 19041 26140
rect 18977 26080 19041 26084
rect 19057 26140 19121 26144
rect 19057 26084 19061 26140
rect 19061 26084 19117 26140
rect 19117 26084 19121 26140
rect 19057 26080 19121 26084
rect 19137 26140 19201 26144
rect 19137 26084 19141 26140
rect 19141 26084 19197 26140
rect 19197 26084 19201 26140
rect 19137 26080 19201 26084
rect 19217 26140 19281 26144
rect 19217 26084 19221 26140
rect 19221 26084 19277 26140
rect 19277 26084 19281 26140
rect 19217 26080 19281 26084
rect 25923 26140 25987 26144
rect 25923 26084 25927 26140
rect 25927 26084 25983 26140
rect 25983 26084 25987 26140
rect 25923 26080 25987 26084
rect 26003 26140 26067 26144
rect 26003 26084 26007 26140
rect 26007 26084 26063 26140
rect 26063 26084 26067 26140
rect 26003 26080 26067 26084
rect 26083 26140 26147 26144
rect 26083 26084 26087 26140
rect 26087 26084 26143 26140
rect 26143 26084 26147 26140
rect 26083 26080 26147 26084
rect 26163 26140 26227 26144
rect 26163 26084 26167 26140
rect 26167 26084 26223 26140
rect 26223 26084 26227 26140
rect 26163 26080 26227 26084
rect 4425 25596 4489 25600
rect 4425 25540 4429 25596
rect 4429 25540 4485 25596
rect 4485 25540 4489 25596
rect 4425 25536 4489 25540
rect 4505 25596 4569 25600
rect 4505 25540 4509 25596
rect 4509 25540 4565 25596
rect 4565 25540 4569 25596
rect 4505 25536 4569 25540
rect 4585 25596 4649 25600
rect 4585 25540 4589 25596
rect 4589 25540 4645 25596
rect 4645 25540 4649 25596
rect 4585 25536 4649 25540
rect 4665 25596 4729 25600
rect 4665 25540 4669 25596
rect 4669 25540 4725 25596
rect 4725 25540 4729 25596
rect 4665 25536 4729 25540
rect 11371 25596 11435 25600
rect 11371 25540 11375 25596
rect 11375 25540 11431 25596
rect 11431 25540 11435 25596
rect 11371 25536 11435 25540
rect 11451 25596 11515 25600
rect 11451 25540 11455 25596
rect 11455 25540 11511 25596
rect 11511 25540 11515 25596
rect 11451 25536 11515 25540
rect 11531 25596 11595 25600
rect 11531 25540 11535 25596
rect 11535 25540 11591 25596
rect 11591 25540 11595 25596
rect 11531 25536 11595 25540
rect 11611 25596 11675 25600
rect 11611 25540 11615 25596
rect 11615 25540 11671 25596
rect 11671 25540 11675 25596
rect 11611 25536 11675 25540
rect 18317 25596 18381 25600
rect 18317 25540 18321 25596
rect 18321 25540 18377 25596
rect 18377 25540 18381 25596
rect 18317 25536 18381 25540
rect 18397 25596 18461 25600
rect 18397 25540 18401 25596
rect 18401 25540 18457 25596
rect 18457 25540 18461 25596
rect 18397 25536 18461 25540
rect 18477 25596 18541 25600
rect 18477 25540 18481 25596
rect 18481 25540 18537 25596
rect 18537 25540 18541 25596
rect 18477 25536 18541 25540
rect 18557 25596 18621 25600
rect 18557 25540 18561 25596
rect 18561 25540 18617 25596
rect 18617 25540 18621 25596
rect 18557 25536 18621 25540
rect 25263 25596 25327 25600
rect 25263 25540 25267 25596
rect 25267 25540 25323 25596
rect 25323 25540 25327 25596
rect 25263 25536 25327 25540
rect 25343 25596 25407 25600
rect 25343 25540 25347 25596
rect 25347 25540 25403 25596
rect 25403 25540 25407 25596
rect 25343 25536 25407 25540
rect 25423 25596 25487 25600
rect 25423 25540 25427 25596
rect 25427 25540 25483 25596
rect 25483 25540 25487 25596
rect 25423 25536 25487 25540
rect 25503 25596 25567 25600
rect 25503 25540 25507 25596
rect 25507 25540 25563 25596
rect 25563 25540 25567 25596
rect 25503 25536 25567 25540
rect 5085 25052 5149 25056
rect 5085 24996 5089 25052
rect 5089 24996 5145 25052
rect 5145 24996 5149 25052
rect 5085 24992 5149 24996
rect 5165 25052 5229 25056
rect 5165 24996 5169 25052
rect 5169 24996 5225 25052
rect 5225 24996 5229 25052
rect 5165 24992 5229 24996
rect 5245 25052 5309 25056
rect 5245 24996 5249 25052
rect 5249 24996 5305 25052
rect 5305 24996 5309 25052
rect 5245 24992 5309 24996
rect 5325 25052 5389 25056
rect 5325 24996 5329 25052
rect 5329 24996 5385 25052
rect 5385 24996 5389 25052
rect 5325 24992 5389 24996
rect 12031 25052 12095 25056
rect 12031 24996 12035 25052
rect 12035 24996 12091 25052
rect 12091 24996 12095 25052
rect 12031 24992 12095 24996
rect 12111 25052 12175 25056
rect 12111 24996 12115 25052
rect 12115 24996 12171 25052
rect 12171 24996 12175 25052
rect 12111 24992 12175 24996
rect 12191 25052 12255 25056
rect 12191 24996 12195 25052
rect 12195 24996 12251 25052
rect 12251 24996 12255 25052
rect 12191 24992 12255 24996
rect 12271 25052 12335 25056
rect 12271 24996 12275 25052
rect 12275 24996 12331 25052
rect 12331 24996 12335 25052
rect 12271 24992 12335 24996
rect 18977 25052 19041 25056
rect 18977 24996 18981 25052
rect 18981 24996 19037 25052
rect 19037 24996 19041 25052
rect 18977 24992 19041 24996
rect 19057 25052 19121 25056
rect 19057 24996 19061 25052
rect 19061 24996 19117 25052
rect 19117 24996 19121 25052
rect 19057 24992 19121 24996
rect 19137 25052 19201 25056
rect 19137 24996 19141 25052
rect 19141 24996 19197 25052
rect 19197 24996 19201 25052
rect 19137 24992 19201 24996
rect 19217 25052 19281 25056
rect 19217 24996 19221 25052
rect 19221 24996 19277 25052
rect 19277 24996 19281 25052
rect 19217 24992 19281 24996
rect 25923 25052 25987 25056
rect 25923 24996 25927 25052
rect 25927 24996 25983 25052
rect 25983 24996 25987 25052
rect 25923 24992 25987 24996
rect 26003 25052 26067 25056
rect 26003 24996 26007 25052
rect 26007 24996 26063 25052
rect 26063 24996 26067 25052
rect 26003 24992 26067 24996
rect 26083 25052 26147 25056
rect 26083 24996 26087 25052
rect 26087 24996 26143 25052
rect 26143 24996 26147 25052
rect 26083 24992 26147 24996
rect 26163 25052 26227 25056
rect 26163 24996 26167 25052
rect 26167 24996 26223 25052
rect 26223 24996 26227 25052
rect 26163 24992 26227 24996
rect 4425 24508 4489 24512
rect 4425 24452 4429 24508
rect 4429 24452 4485 24508
rect 4485 24452 4489 24508
rect 4425 24448 4489 24452
rect 4505 24508 4569 24512
rect 4505 24452 4509 24508
rect 4509 24452 4565 24508
rect 4565 24452 4569 24508
rect 4505 24448 4569 24452
rect 4585 24508 4649 24512
rect 4585 24452 4589 24508
rect 4589 24452 4645 24508
rect 4645 24452 4649 24508
rect 4585 24448 4649 24452
rect 4665 24508 4729 24512
rect 4665 24452 4669 24508
rect 4669 24452 4725 24508
rect 4725 24452 4729 24508
rect 4665 24448 4729 24452
rect 11371 24508 11435 24512
rect 11371 24452 11375 24508
rect 11375 24452 11431 24508
rect 11431 24452 11435 24508
rect 11371 24448 11435 24452
rect 11451 24508 11515 24512
rect 11451 24452 11455 24508
rect 11455 24452 11511 24508
rect 11511 24452 11515 24508
rect 11451 24448 11515 24452
rect 11531 24508 11595 24512
rect 11531 24452 11535 24508
rect 11535 24452 11591 24508
rect 11591 24452 11595 24508
rect 11531 24448 11595 24452
rect 11611 24508 11675 24512
rect 11611 24452 11615 24508
rect 11615 24452 11671 24508
rect 11671 24452 11675 24508
rect 11611 24448 11675 24452
rect 18317 24508 18381 24512
rect 18317 24452 18321 24508
rect 18321 24452 18377 24508
rect 18377 24452 18381 24508
rect 18317 24448 18381 24452
rect 18397 24508 18461 24512
rect 18397 24452 18401 24508
rect 18401 24452 18457 24508
rect 18457 24452 18461 24508
rect 18397 24448 18461 24452
rect 18477 24508 18541 24512
rect 18477 24452 18481 24508
rect 18481 24452 18537 24508
rect 18537 24452 18541 24508
rect 18477 24448 18541 24452
rect 18557 24508 18621 24512
rect 18557 24452 18561 24508
rect 18561 24452 18617 24508
rect 18617 24452 18621 24508
rect 18557 24448 18621 24452
rect 25263 24508 25327 24512
rect 25263 24452 25267 24508
rect 25267 24452 25323 24508
rect 25323 24452 25327 24508
rect 25263 24448 25327 24452
rect 25343 24508 25407 24512
rect 25343 24452 25347 24508
rect 25347 24452 25403 24508
rect 25403 24452 25407 24508
rect 25343 24448 25407 24452
rect 25423 24508 25487 24512
rect 25423 24452 25427 24508
rect 25427 24452 25483 24508
rect 25483 24452 25487 24508
rect 25423 24448 25487 24452
rect 25503 24508 25567 24512
rect 25503 24452 25507 24508
rect 25507 24452 25563 24508
rect 25563 24452 25567 24508
rect 25503 24448 25567 24452
rect 5085 23964 5149 23968
rect 5085 23908 5089 23964
rect 5089 23908 5145 23964
rect 5145 23908 5149 23964
rect 5085 23904 5149 23908
rect 5165 23964 5229 23968
rect 5165 23908 5169 23964
rect 5169 23908 5225 23964
rect 5225 23908 5229 23964
rect 5165 23904 5229 23908
rect 5245 23964 5309 23968
rect 5245 23908 5249 23964
rect 5249 23908 5305 23964
rect 5305 23908 5309 23964
rect 5245 23904 5309 23908
rect 5325 23964 5389 23968
rect 5325 23908 5329 23964
rect 5329 23908 5385 23964
rect 5385 23908 5389 23964
rect 5325 23904 5389 23908
rect 12031 23964 12095 23968
rect 12031 23908 12035 23964
rect 12035 23908 12091 23964
rect 12091 23908 12095 23964
rect 12031 23904 12095 23908
rect 12111 23964 12175 23968
rect 12111 23908 12115 23964
rect 12115 23908 12171 23964
rect 12171 23908 12175 23964
rect 12111 23904 12175 23908
rect 12191 23964 12255 23968
rect 12191 23908 12195 23964
rect 12195 23908 12251 23964
rect 12251 23908 12255 23964
rect 12191 23904 12255 23908
rect 12271 23964 12335 23968
rect 12271 23908 12275 23964
rect 12275 23908 12331 23964
rect 12331 23908 12335 23964
rect 12271 23904 12335 23908
rect 18977 23964 19041 23968
rect 18977 23908 18981 23964
rect 18981 23908 19037 23964
rect 19037 23908 19041 23964
rect 18977 23904 19041 23908
rect 19057 23964 19121 23968
rect 19057 23908 19061 23964
rect 19061 23908 19117 23964
rect 19117 23908 19121 23964
rect 19057 23904 19121 23908
rect 19137 23964 19201 23968
rect 19137 23908 19141 23964
rect 19141 23908 19197 23964
rect 19197 23908 19201 23964
rect 19137 23904 19201 23908
rect 19217 23964 19281 23968
rect 19217 23908 19221 23964
rect 19221 23908 19277 23964
rect 19277 23908 19281 23964
rect 19217 23904 19281 23908
rect 25923 23964 25987 23968
rect 25923 23908 25927 23964
rect 25927 23908 25983 23964
rect 25983 23908 25987 23964
rect 25923 23904 25987 23908
rect 26003 23964 26067 23968
rect 26003 23908 26007 23964
rect 26007 23908 26063 23964
rect 26063 23908 26067 23964
rect 26003 23904 26067 23908
rect 26083 23964 26147 23968
rect 26083 23908 26087 23964
rect 26087 23908 26143 23964
rect 26143 23908 26147 23964
rect 26083 23904 26147 23908
rect 26163 23964 26227 23968
rect 26163 23908 26167 23964
rect 26167 23908 26223 23964
rect 26223 23908 26227 23964
rect 26163 23904 26227 23908
rect 4425 23420 4489 23424
rect 4425 23364 4429 23420
rect 4429 23364 4485 23420
rect 4485 23364 4489 23420
rect 4425 23360 4489 23364
rect 4505 23420 4569 23424
rect 4505 23364 4509 23420
rect 4509 23364 4565 23420
rect 4565 23364 4569 23420
rect 4505 23360 4569 23364
rect 4585 23420 4649 23424
rect 4585 23364 4589 23420
rect 4589 23364 4645 23420
rect 4645 23364 4649 23420
rect 4585 23360 4649 23364
rect 4665 23420 4729 23424
rect 4665 23364 4669 23420
rect 4669 23364 4725 23420
rect 4725 23364 4729 23420
rect 4665 23360 4729 23364
rect 11371 23420 11435 23424
rect 11371 23364 11375 23420
rect 11375 23364 11431 23420
rect 11431 23364 11435 23420
rect 11371 23360 11435 23364
rect 11451 23420 11515 23424
rect 11451 23364 11455 23420
rect 11455 23364 11511 23420
rect 11511 23364 11515 23420
rect 11451 23360 11515 23364
rect 11531 23420 11595 23424
rect 11531 23364 11535 23420
rect 11535 23364 11591 23420
rect 11591 23364 11595 23420
rect 11531 23360 11595 23364
rect 11611 23420 11675 23424
rect 11611 23364 11615 23420
rect 11615 23364 11671 23420
rect 11671 23364 11675 23420
rect 11611 23360 11675 23364
rect 18317 23420 18381 23424
rect 18317 23364 18321 23420
rect 18321 23364 18377 23420
rect 18377 23364 18381 23420
rect 18317 23360 18381 23364
rect 18397 23420 18461 23424
rect 18397 23364 18401 23420
rect 18401 23364 18457 23420
rect 18457 23364 18461 23420
rect 18397 23360 18461 23364
rect 18477 23420 18541 23424
rect 18477 23364 18481 23420
rect 18481 23364 18537 23420
rect 18537 23364 18541 23420
rect 18477 23360 18541 23364
rect 18557 23420 18621 23424
rect 18557 23364 18561 23420
rect 18561 23364 18617 23420
rect 18617 23364 18621 23420
rect 18557 23360 18621 23364
rect 25263 23420 25327 23424
rect 25263 23364 25267 23420
rect 25267 23364 25323 23420
rect 25323 23364 25327 23420
rect 25263 23360 25327 23364
rect 25343 23420 25407 23424
rect 25343 23364 25347 23420
rect 25347 23364 25403 23420
rect 25403 23364 25407 23420
rect 25343 23360 25407 23364
rect 25423 23420 25487 23424
rect 25423 23364 25427 23420
rect 25427 23364 25483 23420
rect 25483 23364 25487 23420
rect 25423 23360 25487 23364
rect 25503 23420 25567 23424
rect 25503 23364 25507 23420
rect 25507 23364 25563 23420
rect 25563 23364 25567 23420
rect 25503 23360 25567 23364
rect 5085 22876 5149 22880
rect 5085 22820 5089 22876
rect 5089 22820 5145 22876
rect 5145 22820 5149 22876
rect 5085 22816 5149 22820
rect 5165 22876 5229 22880
rect 5165 22820 5169 22876
rect 5169 22820 5225 22876
rect 5225 22820 5229 22876
rect 5165 22816 5229 22820
rect 5245 22876 5309 22880
rect 5245 22820 5249 22876
rect 5249 22820 5305 22876
rect 5305 22820 5309 22876
rect 5245 22816 5309 22820
rect 5325 22876 5389 22880
rect 5325 22820 5329 22876
rect 5329 22820 5385 22876
rect 5385 22820 5389 22876
rect 5325 22816 5389 22820
rect 12031 22876 12095 22880
rect 12031 22820 12035 22876
rect 12035 22820 12091 22876
rect 12091 22820 12095 22876
rect 12031 22816 12095 22820
rect 12111 22876 12175 22880
rect 12111 22820 12115 22876
rect 12115 22820 12171 22876
rect 12171 22820 12175 22876
rect 12111 22816 12175 22820
rect 12191 22876 12255 22880
rect 12191 22820 12195 22876
rect 12195 22820 12251 22876
rect 12251 22820 12255 22876
rect 12191 22816 12255 22820
rect 12271 22876 12335 22880
rect 12271 22820 12275 22876
rect 12275 22820 12331 22876
rect 12331 22820 12335 22876
rect 12271 22816 12335 22820
rect 18977 22876 19041 22880
rect 18977 22820 18981 22876
rect 18981 22820 19037 22876
rect 19037 22820 19041 22876
rect 18977 22816 19041 22820
rect 19057 22876 19121 22880
rect 19057 22820 19061 22876
rect 19061 22820 19117 22876
rect 19117 22820 19121 22876
rect 19057 22816 19121 22820
rect 19137 22876 19201 22880
rect 19137 22820 19141 22876
rect 19141 22820 19197 22876
rect 19197 22820 19201 22876
rect 19137 22816 19201 22820
rect 19217 22876 19281 22880
rect 19217 22820 19221 22876
rect 19221 22820 19277 22876
rect 19277 22820 19281 22876
rect 19217 22816 19281 22820
rect 25923 22876 25987 22880
rect 25923 22820 25927 22876
rect 25927 22820 25983 22876
rect 25983 22820 25987 22876
rect 25923 22816 25987 22820
rect 26003 22876 26067 22880
rect 26003 22820 26007 22876
rect 26007 22820 26063 22876
rect 26063 22820 26067 22876
rect 26003 22816 26067 22820
rect 26083 22876 26147 22880
rect 26083 22820 26087 22876
rect 26087 22820 26143 22876
rect 26143 22820 26147 22876
rect 26083 22816 26147 22820
rect 26163 22876 26227 22880
rect 26163 22820 26167 22876
rect 26167 22820 26223 22876
rect 26223 22820 26227 22876
rect 26163 22816 26227 22820
rect 4425 22332 4489 22336
rect 4425 22276 4429 22332
rect 4429 22276 4485 22332
rect 4485 22276 4489 22332
rect 4425 22272 4489 22276
rect 4505 22332 4569 22336
rect 4505 22276 4509 22332
rect 4509 22276 4565 22332
rect 4565 22276 4569 22332
rect 4505 22272 4569 22276
rect 4585 22332 4649 22336
rect 4585 22276 4589 22332
rect 4589 22276 4645 22332
rect 4645 22276 4649 22332
rect 4585 22272 4649 22276
rect 4665 22332 4729 22336
rect 4665 22276 4669 22332
rect 4669 22276 4725 22332
rect 4725 22276 4729 22332
rect 4665 22272 4729 22276
rect 11371 22332 11435 22336
rect 11371 22276 11375 22332
rect 11375 22276 11431 22332
rect 11431 22276 11435 22332
rect 11371 22272 11435 22276
rect 11451 22332 11515 22336
rect 11451 22276 11455 22332
rect 11455 22276 11511 22332
rect 11511 22276 11515 22332
rect 11451 22272 11515 22276
rect 11531 22332 11595 22336
rect 11531 22276 11535 22332
rect 11535 22276 11591 22332
rect 11591 22276 11595 22332
rect 11531 22272 11595 22276
rect 11611 22332 11675 22336
rect 11611 22276 11615 22332
rect 11615 22276 11671 22332
rect 11671 22276 11675 22332
rect 11611 22272 11675 22276
rect 18317 22332 18381 22336
rect 18317 22276 18321 22332
rect 18321 22276 18377 22332
rect 18377 22276 18381 22332
rect 18317 22272 18381 22276
rect 18397 22332 18461 22336
rect 18397 22276 18401 22332
rect 18401 22276 18457 22332
rect 18457 22276 18461 22332
rect 18397 22272 18461 22276
rect 18477 22332 18541 22336
rect 18477 22276 18481 22332
rect 18481 22276 18537 22332
rect 18537 22276 18541 22332
rect 18477 22272 18541 22276
rect 18557 22332 18621 22336
rect 18557 22276 18561 22332
rect 18561 22276 18617 22332
rect 18617 22276 18621 22332
rect 18557 22272 18621 22276
rect 25263 22332 25327 22336
rect 25263 22276 25267 22332
rect 25267 22276 25323 22332
rect 25323 22276 25327 22332
rect 25263 22272 25327 22276
rect 25343 22332 25407 22336
rect 25343 22276 25347 22332
rect 25347 22276 25403 22332
rect 25403 22276 25407 22332
rect 25343 22272 25407 22276
rect 25423 22332 25487 22336
rect 25423 22276 25427 22332
rect 25427 22276 25483 22332
rect 25483 22276 25487 22332
rect 25423 22272 25487 22276
rect 25503 22332 25567 22336
rect 25503 22276 25507 22332
rect 25507 22276 25563 22332
rect 25563 22276 25567 22332
rect 25503 22272 25567 22276
rect 5085 21788 5149 21792
rect 5085 21732 5089 21788
rect 5089 21732 5145 21788
rect 5145 21732 5149 21788
rect 5085 21728 5149 21732
rect 5165 21788 5229 21792
rect 5165 21732 5169 21788
rect 5169 21732 5225 21788
rect 5225 21732 5229 21788
rect 5165 21728 5229 21732
rect 5245 21788 5309 21792
rect 5245 21732 5249 21788
rect 5249 21732 5305 21788
rect 5305 21732 5309 21788
rect 5245 21728 5309 21732
rect 5325 21788 5389 21792
rect 5325 21732 5329 21788
rect 5329 21732 5385 21788
rect 5385 21732 5389 21788
rect 5325 21728 5389 21732
rect 12031 21788 12095 21792
rect 12031 21732 12035 21788
rect 12035 21732 12091 21788
rect 12091 21732 12095 21788
rect 12031 21728 12095 21732
rect 12111 21788 12175 21792
rect 12111 21732 12115 21788
rect 12115 21732 12171 21788
rect 12171 21732 12175 21788
rect 12111 21728 12175 21732
rect 12191 21788 12255 21792
rect 12191 21732 12195 21788
rect 12195 21732 12251 21788
rect 12251 21732 12255 21788
rect 12191 21728 12255 21732
rect 12271 21788 12335 21792
rect 12271 21732 12275 21788
rect 12275 21732 12331 21788
rect 12331 21732 12335 21788
rect 12271 21728 12335 21732
rect 18977 21788 19041 21792
rect 18977 21732 18981 21788
rect 18981 21732 19037 21788
rect 19037 21732 19041 21788
rect 18977 21728 19041 21732
rect 19057 21788 19121 21792
rect 19057 21732 19061 21788
rect 19061 21732 19117 21788
rect 19117 21732 19121 21788
rect 19057 21728 19121 21732
rect 19137 21788 19201 21792
rect 19137 21732 19141 21788
rect 19141 21732 19197 21788
rect 19197 21732 19201 21788
rect 19137 21728 19201 21732
rect 19217 21788 19281 21792
rect 19217 21732 19221 21788
rect 19221 21732 19277 21788
rect 19277 21732 19281 21788
rect 19217 21728 19281 21732
rect 25923 21788 25987 21792
rect 25923 21732 25927 21788
rect 25927 21732 25983 21788
rect 25983 21732 25987 21788
rect 25923 21728 25987 21732
rect 26003 21788 26067 21792
rect 26003 21732 26007 21788
rect 26007 21732 26063 21788
rect 26063 21732 26067 21788
rect 26003 21728 26067 21732
rect 26083 21788 26147 21792
rect 26083 21732 26087 21788
rect 26087 21732 26143 21788
rect 26143 21732 26147 21788
rect 26083 21728 26147 21732
rect 26163 21788 26227 21792
rect 26163 21732 26167 21788
rect 26167 21732 26223 21788
rect 26223 21732 26227 21788
rect 26163 21728 26227 21732
rect 4425 21244 4489 21248
rect 4425 21188 4429 21244
rect 4429 21188 4485 21244
rect 4485 21188 4489 21244
rect 4425 21184 4489 21188
rect 4505 21244 4569 21248
rect 4505 21188 4509 21244
rect 4509 21188 4565 21244
rect 4565 21188 4569 21244
rect 4505 21184 4569 21188
rect 4585 21244 4649 21248
rect 4585 21188 4589 21244
rect 4589 21188 4645 21244
rect 4645 21188 4649 21244
rect 4585 21184 4649 21188
rect 4665 21244 4729 21248
rect 4665 21188 4669 21244
rect 4669 21188 4725 21244
rect 4725 21188 4729 21244
rect 4665 21184 4729 21188
rect 11371 21244 11435 21248
rect 11371 21188 11375 21244
rect 11375 21188 11431 21244
rect 11431 21188 11435 21244
rect 11371 21184 11435 21188
rect 11451 21244 11515 21248
rect 11451 21188 11455 21244
rect 11455 21188 11511 21244
rect 11511 21188 11515 21244
rect 11451 21184 11515 21188
rect 11531 21244 11595 21248
rect 11531 21188 11535 21244
rect 11535 21188 11591 21244
rect 11591 21188 11595 21244
rect 11531 21184 11595 21188
rect 11611 21244 11675 21248
rect 11611 21188 11615 21244
rect 11615 21188 11671 21244
rect 11671 21188 11675 21244
rect 11611 21184 11675 21188
rect 18317 21244 18381 21248
rect 18317 21188 18321 21244
rect 18321 21188 18377 21244
rect 18377 21188 18381 21244
rect 18317 21184 18381 21188
rect 18397 21244 18461 21248
rect 18397 21188 18401 21244
rect 18401 21188 18457 21244
rect 18457 21188 18461 21244
rect 18397 21184 18461 21188
rect 18477 21244 18541 21248
rect 18477 21188 18481 21244
rect 18481 21188 18537 21244
rect 18537 21188 18541 21244
rect 18477 21184 18541 21188
rect 18557 21244 18621 21248
rect 18557 21188 18561 21244
rect 18561 21188 18617 21244
rect 18617 21188 18621 21244
rect 18557 21184 18621 21188
rect 25263 21244 25327 21248
rect 25263 21188 25267 21244
rect 25267 21188 25323 21244
rect 25323 21188 25327 21244
rect 25263 21184 25327 21188
rect 25343 21244 25407 21248
rect 25343 21188 25347 21244
rect 25347 21188 25403 21244
rect 25403 21188 25407 21244
rect 25343 21184 25407 21188
rect 25423 21244 25487 21248
rect 25423 21188 25427 21244
rect 25427 21188 25483 21244
rect 25483 21188 25487 21244
rect 25423 21184 25487 21188
rect 25503 21244 25567 21248
rect 25503 21188 25507 21244
rect 25507 21188 25563 21244
rect 25563 21188 25567 21244
rect 25503 21184 25567 21188
rect 5085 20700 5149 20704
rect 5085 20644 5089 20700
rect 5089 20644 5145 20700
rect 5145 20644 5149 20700
rect 5085 20640 5149 20644
rect 5165 20700 5229 20704
rect 5165 20644 5169 20700
rect 5169 20644 5225 20700
rect 5225 20644 5229 20700
rect 5165 20640 5229 20644
rect 5245 20700 5309 20704
rect 5245 20644 5249 20700
rect 5249 20644 5305 20700
rect 5305 20644 5309 20700
rect 5245 20640 5309 20644
rect 5325 20700 5389 20704
rect 5325 20644 5329 20700
rect 5329 20644 5385 20700
rect 5385 20644 5389 20700
rect 5325 20640 5389 20644
rect 12031 20700 12095 20704
rect 12031 20644 12035 20700
rect 12035 20644 12091 20700
rect 12091 20644 12095 20700
rect 12031 20640 12095 20644
rect 12111 20700 12175 20704
rect 12111 20644 12115 20700
rect 12115 20644 12171 20700
rect 12171 20644 12175 20700
rect 12111 20640 12175 20644
rect 12191 20700 12255 20704
rect 12191 20644 12195 20700
rect 12195 20644 12251 20700
rect 12251 20644 12255 20700
rect 12191 20640 12255 20644
rect 12271 20700 12335 20704
rect 12271 20644 12275 20700
rect 12275 20644 12331 20700
rect 12331 20644 12335 20700
rect 12271 20640 12335 20644
rect 18977 20700 19041 20704
rect 18977 20644 18981 20700
rect 18981 20644 19037 20700
rect 19037 20644 19041 20700
rect 18977 20640 19041 20644
rect 19057 20700 19121 20704
rect 19057 20644 19061 20700
rect 19061 20644 19117 20700
rect 19117 20644 19121 20700
rect 19057 20640 19121 20644
rect 19137 20700 19201 20704
rect 19137 20644 19141 20700
rect 19141 20644 19197 20700
rect 19197 20644 19201 20700
rect 19137 20640 19201 20644
rect 19217 20700 19281 20704
rect 19217 20644 19221 20700
rect 19221 20644 19277 20700
rect 19277 20644 19281 20700
rect 19217 20640 19281 20644
rect 25923 20700 25987 20704
rect 25923 20644 25927 20700
rect 25927 20644 25983 20700
rect 25983 20644 25987 20700
rect 25923 20640 25987 20644
rect 26003 20700 26067 20704
rect 26003 20644 26007 20700
rect 26007 20644 26063 20700
rect 26063 20644 26067 20700
rect 26003 20640 26067 20644
rect 26083 20700 26147 20704
rect 26083 20644 26087 20700
rect 26087 20644 26143 20700
rect 26143 20644 26147 20700
rect 26083 20640 26147 20644
rect 26163 20700 26227 20704
rect 26163 20644 26167 20700
rect 26167 20644 26223 20700
rect 26223 20644 26227 20700
rect 26163 20640 26227 20644
rect 4425 20156 4489 20160
rect 4425 20100 4429 20156
rect 4429 20100 4485 20156
rect 4485 20100 4489 20156
rect 4425 20096 4489 20100
rect 4505 20156 4569 20160
rect 4505 20100 4509 20156
rect 4509 20100 4565 20156
rect 4565 20100 4569 20156
rect 4505 20096 4569 20100
rect 4585 20156 4649 20160
rect 4585 20100 4589 20156
rect 4589 20100 4645 20156
rect 4645 20100 4649 20156
rect 4585 20096 4649 20100
rect 4665 20156 4729 20160
rect 4665 20100 4669 20156
rect 4669 20100 4725 20156
rect 4725 20100 4729 20156
rect 4665 20096 4729 20100
rect 11371 20156 11435 20160
rect 11371 20100 11375 20156
rect 11375 20100 11431 20156
rect 11431 20100 11435 20156
rect 11371 20096 11435 20100
rect 11451 20156 11515 20160
rect 11451 20100 11455 20156
rect 11455 20100 11511 20156
rect 11511 20100 11515 20156
rect 11451 20096 11515 20100
rect 11531 20156 11595 20160
rect 11531 20100 11535 20156
rect 11535 20100 11591 20156
rect 11591 20100 11595 20156
rect 11531 20096 11595 20100
rect 11611 20156 11675 20160
rect 11611 20100 11615 20156
rect 11615 20100 11671 20156
rect 11671 20100 11675 20156
rect 11611 20096 11675 20100
rect 18317 20156 18381 20160
rect 18317 20100 18321 20156
rect 18321 20100 18377 20156
rect 18377 20100 18381 20156
rect 18317 20096 18381 20100
rect 18397 20156 18461 20160
rect 18397 20100 18401 20156
rect 18401 20100 18457 20156
rect 18457 20100 18461 20156
rect 18397 20096 18461 20100
rect 18477 20156 18541 20160
rect 18477 20100 18481 20156
rect 18481 20100 18537 20156
rect 18537 20100 18541 20156
rect 18477 20096 18541 20100
rect 18557 20156 18621 20160
rect 18557 20100 18561 20156
rect 18561 20100 18617 20156
rect 18617 20100 18621 20156
rect 18557 20096 18621 20100
rect 25263 20156 25327 20160
rect 25263 20100 25267 20156
rect 25267 20100 25323 20156
rect 25323 20100 25327 20156
rect 25263 20096 25327 20100
rect 25343 20156 25407 20160
rect 25343 20100 25347 20156
rect 25347 20100 25403 20156
rect 25403 20100 25407 20156
rect 25343 20096 25407 20100
rect 25423 20156 25487 20160
rect 25423 20100 25427 20156
rect 25427 20100 25483 20156
rect 25483 20100 25487 20156
rect 25423 20096 25487 20100
rect 25503 20156 25567 20160
rect 25503 20100 25507 20156
rect 25507 20100 25563 20156
rect 25563 20100 25567 20156
rect 25503 20096 25567 20100
rect 5085 19612 5149 19616
rect 5085 19556 5089 19612
rect 5089 19556 5145 19612
rect 5145 19556 5149 19612
rect 5085 19552 5149 19556
rect 5165 19612 5229 19616
rect 5165 19556 5169 19612
rect 5169 19556 5225 19612
rect 5225 19556 5229 19612
rect 5165 19552 5229 19556
rect 5245 19612 5309 19616
rect 5245 19556 5249 19612
rect 5249 19556 5305 19612
rect 5305 19556 5309 19612
rect 5245 19552 5309 19556
rect 5325 19612 5389 19616
rect 5325 19556 5329 19612
rect 5329 19556 5385 19612
rect 5385 19556 5389 19612
rect 5325 19552 5389 19556
rect 12031 19612 12095 19616
rect 12031 19556 12035 19612
rect 12035 19556 12091 19612
rect 12091 19556 12095 19612
rect 12031 19552 12095 19556
rect 12111 19612 12175 19616
rect 12111 19556 12115 19612
rect 12115 19556 12171 19612
rect 12171 19556 12175 19612
rect 12111 19552 12175 19556
rect 12191 19612 12255 19616
rect 12191 19556 12195 19612
rect 12195 19556 12251 19612
rect 12251 19556 12255 19612
rect 12191 19552 12255 19556
rect 12271 19612 12335 19616
rect 12271 19556 12275 19612
rect 12275 19556 12331 19612
rect 12331 19556 12335 19612
rect 12271 19552 12335 19556
rect 18977 19612 19041 19616
rect 18977 19556 18981 19612
rect 18981 19556 19037 19612
rect 19037 19556 19041 19612
rect 18977 19552 19041 19556
rect 19057 19612 19121 19616
rect 19057 19556 19061 19612
rect 19061 19556 19117 19612
rect 19117 19556 19121 19612
rect 19057 19552 19121 19556
rect 19137 19612 19201 19616
rect 19137 19556 19141 19612
rect 19141 19556 19197 19612
rect 19197 19556 19201 19612
rect 19137 19552 19201 19556
rect 19217 19612 19281 19616
rect 19217 19556 19221 19612
rect 19221 19556 19277 19612
rect 19277 19556 19281 19612
rect 19217 19552 19281 19556
rect 25923 19612 25987 19616
rect 25923 19556 25927 19612
rect 25927 19556 25983 19612
rect 25983 19556 25987 19612
rect 25923 19552 25987 19556
rect 26003 19612 26067 19616
rect 26003 19556 26007 19612
rect 26007 19556 26063 19612
rect 26063 19556 26067 19612
rect 26003 19552 26067 19556
rect 26083 19612 26147 19616
rect 26083 19556 26087 19612
rect 26087 19556 26143 19612
rect 26143 19556 26147 19612
rect 26083 19552 26147 19556
rect 26163 19612 26227 19616
rect 26163 19556 26167 19612
rect 26167 19556 26223 19612
rect 26223 19556 26227 19612
rect 26163 19552 26227 19556
rect 4425 19068 4489 19072
rect 4425 19012 4429 19068
rect 4429 19012 4485 19068
rect 4485 19012 4489 19068
rect 4425 19008 4489 19012
rect 4505 19068 4569 19072
rect 4505 19012 4509 19068
rect 4509 19012 4565 19068
rect 4565 19012 4569 19068
rect 4505 19008 4569 19012
rect 4585 19068 4649 19072
rect 4585 19012 4589 19068
rect 4589 19012 4645 19068
rect 4645 19012 4649 19068
rect 4585 19008 4649 19012
rect 4665 19068 4729 19072
rect 4665 19012 4669 19068
rect 4669 19012 4725 19068
rect 4725 19012 4729 19068
rect 4665 19008 4729 19012
rect 11371 19068 11435 19072
rect 11371 19012 11375 19068
rect 11375 19012 11431 19068
rect 11431 19012 11435 19068
rect 11371 19008 11435 19012
rect 11451 19068 11515 19072
rect 11451 19012 11455 19068
rect 11455 19012 11511 19068
rect 11511 19012 11515 19068
rect 11451 19008 11515 19012
rect 11531 19068 11595 19072
rect 11531 19012 11535 19068
rect 11535 19012 11591 19068
rect 11591 19012 11595 19068
rect 11531 19008 11595 19012
rect 11611 19068 11675 19072
rect 11611 19012 11615 19068
rect 11615 19012 11671 19068
rect 11671 19012 11675 19068
rect 11611 19008 11675 19012
rect 18317 19068 18381 19072
rect 18317 19012 18321 19068
rect 18321 19012 18377 19068
rect 18377 19012 18381 19068
rect 18317 19008 18381 19012
rect 18397 19068 18461 19072
rect 18397 19012 18401 19068
rect 18401 19012 18457 19068
rect 18457 19012 18461 19068
rect 18397 19008 18461 19012
rect 18477 19068 18541 19072
rect 18477 19012 18481 19068
rect 18481 19012 18537 19068
rect 18537 19012 18541 19068
rect 18477 19008 18541 19012
rect 18557 19068 18621 19072
rect 18557 19012 18561 19068
rect 18561 19012 18617 19068
rect 18617 19012 18621 19068
rect 18557 19008 18621 19012
rect 25263 19068 25327 19072
rect 25263 19012 25267 19068
rect 25267 19012 25323 19068
rect 25323 19012 25327 19068
rect 25263 19008 25327 19012
rect 25343 19068 25407 19072
rect 25343 19012 25347 19068
rect 25347 19012 25403 19068
rect 25403 19012 25407 19068
rect 25343 19008 25407 19012
rect 25423 19068 25487 19072
rect 25423 19012 25427 19068
rect 25427 19012 25483 19068
rect 25483 19012 25487 19068
rect 25423 19008 25487 19012
rect 25503 19068 25567 19072
rect 25503 19012 25507 19068
rect 25507 19012 25563 19068
rect 25563 19012 25567 19068
rect 25503 19008 25567 19012
rect 5085 18524 5149 18528
rect 5085 18468 5089 18524
rect 5089 18468 5145 18524
rect 5145 18468 5149 18524
rect 5085 18464 5149 18468
rect 5165 18524 5229 18528
rect 5165 18468 5169 18524
rect 5169 18468 5225 18524
rect 5225 18468 5229 18524
rect 5165 18464 5229 18468
rect 5245 18524 5309 18528
rect 5245 18468 5249 18524
rect 5249 18468 5305 18524
rect 5305 18468 5309 18524
rect 5245 18464 5309 18468
rect 5325 18524 5389 18528
rect 5325 18468 5329 18524
rect 5329 18468 5385 18524
rect 5385 18468 5389 18524
rect 5325 18464 5389 18468
rect 12031 18524 12095 18528
rect 12031 18468 12035 18524
rect 12035 18468 12091 18524
rect 12091 18468 12095 18524
rect 12031 18464 12095 18468
rect 12111 18524 12175 18528
rect 12111 18468 12115 18524
rect 12115 18468 12171 18524
rect 12171 18468 12175 18524
rect 12111 18464 12175 18468
rect 12191 18524 12255 18528
rect 12191 18468 12195 18524
rect 12195 18468 12251 18524
rect 12251 18468 12255 18524
rect 12191 18464 12255 18468
rect 12271 18524 12335 18528
rect 12271 18468 12275 18524
rect 12275 18468 12331 18524
rect 12331 18468 12335 18524
rect 12271 18464 12335 18468
rect 18977 18524 19041 18528
rect 18977 18468 18981 18524
rect 18981 18468 19037 18524
rect 19037 18468 19041 18524
rect 18977 18464 19041 18468
rect 19057 18524 19121 18528
rect 19057 18468 19061 18524
rect 19061 18468 19117 18524
rect 19117 18468 19121 18524
rect 19057 18464 19121 18468
rect 19137 18524 19201 18528
rect 19137 18468 19141 18524
rect 19141 18468 19197 18524
rect 19197 18468 19201 18524
rect 19137 18464 19201 18468
rect 19217 18524 19281 18528
rect 19217 18468 19221 18524
rect 19221 18468 19277 18524
rect 19277 18468 19281 18524
rect 19217 18464 19281 18468
rect 25923 18524 25987 18528
rect 25923 18468 25927 18524
rect 25927 18468 25983 18524
rect 25983 18468 25987 18524
rect 25923 18464 25987 18468
rect 26003 18524 26067 18528
rect 26003 18468 26007 18524
rect 26007 18468 26063 18524
rect 26063 18468 26067 18524
rect 26003 18464 26067 18468
rect 26083 18524 26147 18528
rect 26083 18468 26087 18524
rect 26087 18468 26143 18524
rect 26143 18468 26147 18524
rect 26083 18464 26147 18468
rect 26163 18524 26227 18528
rect 26163 18468 26167 18524
rect 26167 18468 26223 18524
rect 26223 18468 26227 18524
rect 26163 18464 26227 18468
rect 4425 17980 4489 17984
rect 4425 17924 4429 17980
rect 4429 17924 4485 17980
rect 4485 17924 4489 17980
rect 4425 17920 4489 17924
rect 4505 17980 4569 17984
rect 4505 17924 4509 17980
rect 4509 17924 4565 17980
rect 4565 17924 4569 17980
rect 4505 17920 4569 17924
rect 4585 17980 4649 17984
rect 4585 17924 4589 17980
rect 4589 17924 4645 17980
rect 4645 17924 4649 17980
rect 4585 17920 4649 17924
rect 4665 17980 4729 17984
rect 4665 17924 4669 17980
rect 4669 17924 4725 17980
rect 4725 17924 4729 17980
rect 4665 17920 4729 17924
rect 11371 17980 11435 17984
rect 11371 17924 11375 17980
rect 11375 17924 11431 17980
rect 11431 17924 11435 17980
rect 11371 17920 11435 17924
rect 11451 17980 11515 17984
rect 11451 17924 11455 17980
rect 11455 17924 11511 17980
rect 11511 17924 11515 17980
rect 11451 17920 11515 17924
rect 11531 17980 11595 17984
rect 11531 17924 11535 17980
rect 11535 17924 11591 17980
rect 11591 17924 11595 17980
rect 11531 17920 11595 17924
rect 11611 17980 11675 17984
rect 11611 17924 11615 17980
rect 11615 17924 11671 17980
rect 11671 17924 11675 17980
rect 11611 17920 11675 17924
rect 18317 17980 18381 17984
rect 18317 17924 18321 17980
rect 18321 17924 18377 17980
rect 18377 17924 18381 17980
rect 18317 17920 18381 17924
rect 18397 17980 18461 17984
rect 18397 17924 18401 17980
rect 18401 17924 18457 17980
rect 18457 17924 18461 17980
rect 18397 17920 18461 17924
rect 18477 17980 18541 17984
rect 18477 17924 18481 17980
rect 18481 17924 18537 17980
rect 18537 17924 18541 17980
rect 18477 17920 18541 17924
rect 18557 17980 18621 17984
rect 18557 17924 18561 17980
rect 18561 17924 18617 17980
rect 18617 17924 18621 17980
rect 18557 17920 18621 17924
rect 25263 17980 25327 17984
rect 25263 17924 25267 17980
rect 25267 17924 25323 17980
rect 25323 17924 25327 17980
rect 25263 17920 25327 17924
rect 25343 17980 25407 17984
rect 25343 17924 25347 17980
rect 25347 17924 25403 17980
rect 25403 17924 25407 17980
rect 25343 17920 25407 17924
rect 25423 17980 25487 17984
rect 25423 17924 25427 17980
rect 25427 17924 25483 17980
rect 25483 17924 25487 17980
rect 25423 17920 25487 17924
rect 25503 17980 25567 17984
rect 25503 17924 25507 17980
rect 25507 17924 25563 17980
rect 25563 17924 25567 17980
rect 25503 17920 25567 17924
rect 5085 17436 5149 17440
rect 5085 17380 5089 17436
rect 5089 17380 5145 17436
rect 5145 17380 5149 17436
rect 5085 17376 5149 17380
rect 5165 17436 5229 17440
rect 5165 17380 5169 17436
rect 5169 17380 5225 17436
rect 5225 17380 5229 17436
rect 5165 17376 5229 17380
rect 5245 17436 5309 17440
rect 5245 17380 5249 17436
rect 5249 17380 5305 17436
rect 5305 17380 5309 17436
rect 5245 17376 5309 17380
rect 5325 17436 5389 17440
rect 5325 17380 5329 17436
rect 5329 17380 5385 17436
rect 5385 17380 5389 17436
rect 5325 17376 5389 17380
rect 12031 17436 12095 17440
rect 12031 17380 12035 17436
rect 12035 17380 12091 17436
rect 12091 17380 12095 17436
rect 12031 17376 12095 17380
rect 12111 17436 12175 17440
rect 12111 17380 12115 17436
rect 12115 17380 12171 17436
rect 12171 17380 12175 17436
rect 12111 17376 12175 17380
rect 12191 17436 12255 17440
rect 12191 17380 12195 17436
rect 12195 17380 12251 17436
rect 12251 17380 12255 17436
rect 12191 17376 12255 17380
rect 12271 17436 12335 17440
rect 12271 17380 12275 17436
rect 12275 17380 12331 17436
rect 12331 17380 12335 17436
rect 12271 17376 12335 17380
rect 18977 17436 19041 17440
rect 18977 17380 18981 17436
rect 18981 17380 19037 17436
rect 19037 17380 19041 17436
rect 18977 17376 19041 17380
rect 19057 17436 19121 17440
rect 19057 17380 19061 17436
rect 19061 17380 19117 17436
rect 19117 17380 19121 17436
rect 19057 17376 19121 17380
rect 19137 17436 19201 17440
rect 19137 17380 19141 17436
rect 19141 17380 19197 17436
rect 19197 17380 19201 17436
rect 19137 17376 19201 17380
rect 19217 17436 19281 17440
rect 19217 17380 19221 17436
rect 19221 17380 19277 17436
rect 19277 17380 19281 17436
rect 19217 17376 19281 17380
rect 25923 17436 25987 17440
rect 25923 17380 25927 17436
rect 25927 17380 25983 17436
rect 25983 17380 25987 17436
rect 25923 17376 25987 17380
rect 26003 17436 26067 17440
rect 26003 17380 26007 17436
rect 26007 17380 26063 17436
rect 26063 17380 26067 17436
rect 26003 17376 26067 17380
rect 26083 17436 26147 17440
rect 26083 17380 26087 17436
rect 26087 17380 26143 17436
rect 26143 17380 26147 17436
rect 26083 17376 26147 17380
rect 26163 17436 26227 17440
rect 26163 17380 26167 17436
rect 26167 17380 26223 17436
rect 26223 17380 26227 17436
rect 26163 17376 26227 17380
rect 4425 16892 4489 16896
rect 4425 16836 4429 16892
rect 4429 16836 4485 16892
rect 4485 16836 4489 16892
rect 4425 16832 4489 16836
rect 4505 16892 4569 16896
rect 4505 16836 4509 16892
rect 4509 16836 4565 16892
rect 4565 16836 4569 16892
rect 4505 16832 4569 16836
rect 4585 16892 4649 16896
rect 4585 16836 4589 16892
rect 4589 16836 4645 16892
rect 4645 16836 4649 16892
rect 4585 16832 4649 16836
rect 4665 16892 4729 16896
rect 4665 16836 4669 16892
rect 4669 16836 4725 16892
rect 4725 16836 4729 16892
rect 4665 16832 4729 16836
rect 11371 16892 11435 16896
rect 11371 16836 11375 16892
rect 11375 16836 11431 16892
rect 11431 16836 11435 16892
rect 11371 16832 11435 16836
rect 11451 16892 11515 16896
rect 11451 16836 11455 16892
rect 11455 16836 11511 16892
rect 11511 16836 11515 16892
rect 11451 16832 11515 16836
rect 11531 16892 11595 16896
rect 11531 16836 11535 16892
rect 11535 16836 11591 16892
rect 11591 16836 11595 16892
rect 11531 16832 11595 16836
rect 11611 16892 11675 16896
rect 11611 16836 11615 16892
rect 11615 16836 11671 16892
rect 11671 16836 11675 16892
rect 11611 16832 11675 16836
rect 18317 16892 18381 16896
rect 18317 16836 18321 16892
rect 18321 16836 18377 16892
rect 18377 16836 18381 16892
rect 18317 16832 18381 16836
rect 18397 16892 18461 16896
rect 18397 16836 18401 16892
rect 18401 16836 18457 16892
rect 18457 16836 18461 16892
rect 18397 16832 18461 16836
rect 18477 16892 18541 16896
rect 18477 16836 18481 16892
rect 18481 16836 18537 16892
rect 18537 16836 18541 16892
rect 18477 16832 18541 16836
rect 18557 16892 18621 16896
rect 18557 16836 18561 16892
rect 18561 16836 18617 16892
rect 18617 16836 18621 16892
rect 18557 16832 18621 16836
rect 25263 16892 25327 16896
rect 25263 16836 25267 16892
rect 25267 16836 25323 16892
rect 25323 16836 25327 16892
rect 25263 16832 25327 16836
rect 25343 16892 25407 16896
rect 25343 16836 25347 16892
rect 25347 16836 25403 16892
rect 25403 16836 25407 16892
rect 25343 16832 25407 16836
rect 25423 16892 25487 16896
rect 25423 16836 25427 16892
rect 25427 16836 25483 16892
rect 25483 16836 25487 16892
rect 25423 16832 25487 16836
rect 25503 16892 25567 16896
rect 25503 16836 25507 16892
rect 25507 16836 25563 16892
rect 25563 16836 25567 16892
rect 25503 16832 25567 16836
rect 5085 16348 5149 16352
rect 5085 16292 5089 16348
rect 5089 16292 5145 16348
rect 5145 16292 5149 16348
rect 5085 16288 5149 16292
rect 5165 16348 5229 16352
rect 5165 16292 5169 16348
rect 5169 16292 5225 16348
rect 5225 16292 5229 16348
rect 5165 16288 5229 16292
rect 5245 16348 5309 16352
rect 5245 16292 5249 16348
rect 5249 16292 5305 16348
rect 5305 16292 5309 16348
rect 5245 16288 5309 16292
rect 5325 16348 5389 16352
rect 5325 16292 5329 16348
rect 5329 16292 5385 16348
rect 5385 16292 5389 16348
rect 5325 16288 5389 16292
rect 12031 16348 12095 16352
rect 12031 16292 12035 16348
rect 12035 16292 12091 16348
rect 12091 16292 12095 16348
rect 12031 16288 12095 16292
rect 12111 16348 12175 16352
rect 12111 16292 12115 16348
rect 12115 16292 12171 16348
rect 12171 16292 12175 16348
rect 12111 16288 12175 16292
rect 12191 16348 12255 16352
rect 12191 16292 12195 16348
rect 12195 16292 12251 16348
rect 12251 16292 12255 16348
rect 12191 16288 12255 16292
rect 12271 16348 12335 16352
rect 12271 16292 12275 16348
rect 12275 16292 12331 16348
rect 12331 16292 12335 16348
rect 12271 16288 12335 16292
rect 18977 16348 19041 16352
rect 18977 16292 18981 16348
rect 18981 16292 19037 16348
rect 19037 16292 19041 16348
rect 18977 16288 19041 16292
rect 19057 16348 19121 16352
rect 19057 16292 19061 16348
rect 19061 16292 19117 16348
rect 19117 16292 19121 16348
rect 19057 16288 19121 16292
rect 19137 16348 19201 16352
rect 19137 16292 19141 16348
rect 19141 16292 19197 16348
rect 19197 16292 19201 16348
rect 19137 16288 19201 16292
rect 19217 16348 19281 16352
rect 19217 16292 19221 16348
rect 19221 16292 19277 16348
rect 19277 16292 19281 16348
rect 19217 16288 19281 16292
rect 25923 16348 25987 16352
rect 25923 16292 25927 16348
rect 25927 16292 25983 16348
rect 25983 16292 25987 16348
rect 25923 16288 25987 16292
rect 26003 16348 26067 16352
rect 26003 16292 26007 16348
rect 26007 16292 26063 16348
rect 26063 16292 26067 16348
rect 26003 16288 26067 16292
rect 26083 16348 26147 16352
rect 26083 16292 26087 16348
rect 26087 16292 26143 16348
rect 26143 16292 26147 16348
rect 26083 16288 26147 16292
rect 26163 16348 26227 16352
rect 26163 16292 26167 16348
rect 26167 16292 26223 16348
rect 26223 16292 26227 16348
rect 26163 16288 26227 16292
rect 4425 15804 4489 15808
rect 4425 15748 4429 15804
rect 4429 15748 4485 15804
rect 4485 15748 4489 15804
rect 4425 15744 4489 15748
rect 4505 15804 4569 15808
rect 4505 15748 4509 15804
rect 4509 15748 4565 15804
rect 4565 15748 4569 15804
rect 4505 15744 4569 15748
rect 4585 15804 4649 15808
rect 4585 15748 4589 15804
rect 4589 15748 4645 15804
rect 4645 15748 4649 15804
rect 4585 15744 4649 15748
rect 4665 15804 4729 15808
rect 4665 15748 4669 15804
rect 4669 15748 4725 15804
rect 4725 15748 4729 15804
rect 4665 15744 4729 15748
rect 11371 15804 11435 15808
rect 11371 15748 11375 15804
rect 11375 15748 11431 15804
rect 11431 15748 11435 15804
rect 11371 15744 11435 15748
rect 11451 15804 11515 15808
rect 11451 15748 11455 15804
rect 11455 15748 11511 15804
rect 11511 15748 11515 15804
rect 11451 15744 11515 15748
rect 11531 15804 11595 15808
rect 11531 15748 11535 15804
rect 11535 15748 11591 15804
rect 11591 15748 11595 15804
rect 11531 15744 11595 15748
rect 11611 15804 11675 15808
rect 11611 15748 11615 15804
rect 11615 15748 11671 15804
rect 11671 15748 11675 15804
rect 11611 15744 11675 15748
rect 18317 15804 18381 15808
rect 18317 15748 18321 15804
rect 18321 15748 18377 15804
rect 18377 15748 18381 15804
rect 18317 15744 18381 15748
rect 18397 15804 18461 15808
rect 18397 15748 18401 15804
rect 18401 15748 18457 15804
rect 18457 15748 18461 15804
rect 18397 15744 18461 15748
rect 18477 15804 18541 15808
rect 18477 15748 18481 15804
rect 18481 15748 18537 15804
rect 18537 15748 18541 15804
rect 18477 15744 18541 15748
rect 18557 15804 18621 15808
rect 18557 15748 18561 15804
rect 18561 15748 18617 15804
rect 18617 15748 18621 15804
rect 18557 15744 18621 15748
rect 25263 15804 25327 15808
rect 25263 15748 25267 15804
rect 25267 15748 25323 15804
rect 25323 15748 25327 15804
rect 25263 15744 25327 15748
rect 25343 15804 25407 15808
rect 25343 15748 25347 15804
rect 25347 15748 25403 15804
rect 25403 15748 25407 15804
rect 25343 15744 25407 15748
rect 25423 15804 25487 15808
rect 25423 15748 25427 15804
rect 25427 15748 25483 15804
rect 25483 15748 25487 15804
rect 25423 15744 25487 15748
rect 25503 15804 25567 15808
rect 25503 15748 25507 15804
rect 25507 15748 25563 15804
rect 25563 15748 25567 15804
rect 25503 15744 25567 15748
rect 24900 15676 24964 15740
rect 5085 15260 5149 15264
rect 5085 15204 5089 15260
rect 5089 15204 5145 15260
rect 5145 15204 5149 15260
rect 5085 15200 5149 15204
rect 5165 15260 5229 15264
rect 5165 15204 5169 15260
rect 5169 15204 5225 15260
rect 5225 15204 5229 15260
rect 5165 15200 5229 15204
rect 5245 15260 5309 15264
rect 5245 15204 5249 15260
rect 5249 15204 5305 15260
rect 5305 15204 5309 15260
rect 5245 15200 5309 15204
rect 5325 15260 5389 15264
rect 5325 15204 5329 15260
rect 5329 15204 5385 15260
rect 5385 15204 5389 15260
rect 5325 15200 5389 15204
rect 12031 15260 12095 15264
rect 12031 15204 12035 15260
rect 12035 15204 12091 15260
rect 12091 15204 12095 15260
rect 12031 15200 12095 15204
rect 12111 15260 12175 15264
rect 12111 15204 12115 15260
rect 12115 15204 12171 15260
rect 12171 15204 12175 15260
rect 12111 15200 12175 15204
rect 12191 15260 12255 15264
rect 12191 15204 12195 15260
rect 12195 15204 12251 15260
rect 12251 15204 12255 15260
rect 12191 15200 12255 15204
rect 12271 15260 12335 15264
rect 12271 15204 12275 15260
rect 12275 15204 12331 15260
rect 12331 15204 12335 15260
rect 12271 15200 12335 15204
rect 18977 15260 19041 15264
rect 18977 15204 18981 15260
rect 18981 15204 19037 15260
rect 19037 15204 19041 15260
rect 18977 15200 19041 15204
rect 19057 15260 19121 15264
rect 19057 15204 19061 15260
rect 19061 15204 19117 15260
rect 19117 15204 19121 15260
rect 19057 15200 19121 15204
rect 19137 15260 19201 15264
rect 19137 15204 19141 15260
rect 19141 15204 19197 15260
rect 19197 15204 19201 15260
rect 19137 15200 19201 15204
rect 19217 15260 19281 15264
rect 19217 15204 19221 15260
rect 19221 15204 19277 15260
rect 19277 15204 19281 15260
rect 19217 15200 19281 15204
rect 25923 15260 25987 15264
rect 25923 15204 25927 15260
rect 25927 15204 25983 15260
rect 25983 15204 25987 15260
rect 25923 15200 25987 15204
rect 26003 15260 26067 15264
rect 26003 15204 26007 15260
rect 26007 15204 26063 15260
rect 26063 15204 26067 15260
rect 26003 15200 26067 15204
rect 26083 15260 26147 15264
rect 26083 15204 26087 15260
rect 26087 15204 26143 15260
rect 26143 15204 26147 15260
rect 26083 15200 26147 15204
rect 26163 15260 26227 15264
rect 26163 15204 26167 15260
rect 26167 15204 26223 15260
rect 26223 15204 26227 15260
rect 26163 15200 26227 15204
rect 4425 14716 4489 14720
rect 4425 14660 4429 14716
rect 4429 14660 4485 14716
rect 4485 14660 4489 14716
rect 4425 14656 4489 14660
rect 4505 14716 4569 14720
rect 4505 14660 4509 14716
rect 4509 14660 4565 14716
rect 4565 14660 4569 14716
rect 4505 14656 4569 14660
rect 4585 14716 4649 14720
rect 4585 14660 4589 14716
rect 4589 14660 4645 14716
rect 4645 14660 4649 14716
rect 4585 14656 4649 14660
rect 4665 14716 4729 14720
rect 4665 14660 4669 14716
rect 4669 14660 4725 14716
rect 4725 14660 4729 14716
rect 4665 14656 4729 14660
rect 11371 14716 11435 14720
rect 11371 14660 11375 14716
rect 11375 14660 11431 14716
rect 11431 14660 11435 14716
rect 11371 14656 11435 14660
rect 11451 14716 11515 14720
rect 11451 14660 11455 14716
rect 11455 14660 11511 14716
rect 11511 14660 11515 14716
rect 11451 14656 11515 14660
rect 11531 14716 11595 14720
rect 11531 14660 11535 14716
rect 11535 14660 11591 14716
rect 11591 14660 11595 14716
rect 11531 14656 11595 14660
rect 11611 14716 11675 14720
rect 11611 14660 11615 14716
rect 11615 14660 11671 14716
rect 11671 14660 11675 14716
rect 11611 14656 11675 14660
rect 18317 14716 18381 14720
rect 18317 14660 18321 14716
rect 18321 14660 18377 14716
rect 18377 14660 18381 14716
rect 18317 14656 18381 14660
rect 18397 14716 18461 14720
rect 18397 14660 18401 14716
rect 18401 14660 18457 14716
rect 18457 14660 18461 14716
rect 18397 14656 18461 14660
rect 18477 14716 18541 14720
rect 18477 14660 18481 14716
rect 18481 14660 18537 14716
rect 18537 14660 18541 14716
rect 18477 14656 18541 14660
rect 18557 14716 18621 14720
rect 18557 14660 18561 14716
rect 18561 14660 18617 14716
rect 18617 14660 18621 14716
rect 18557 14656 18621 14660
rect 25263 14716 25327 14720
rect 25263 14660 25267 14716
rect 25267 14660 25323 14716
rect 25323 14660 25327 14716
rect 25263 14656 25327 14660
rect 25343 14716 25407 14720
rect 25343 14660 25347 14716
rect 25347 14660 25403 14716
rect 25403 14660 25407 14716
rect 25343 14656 25407 14660
rect 25423 14716 25487 14720
rect 25423 14660 25427 14716
rect 25427 14660 25483 14716
rect 25483 14660 25487 14716
rect 25423 14656 25487 14660
rect 25503 14716 25567 14720
rect 25503 14660 25507 14716
rect 25507 14660 25563 14716
rect 25563 14660 25567 14716
rect 25503 14656 25567 14660
rect 5085 14172 5149 14176
rect 5085 14116 5089 14172
rect 5089 14116 5145 14172
rect 5145 14116 5149 14172
rect 5085 14112 5149 14116
rect 5165 14172 5229 14176
rect 5165 14116 5169 14172
rect 5169 14116 5225 14172
rect 5225 14116 5229 14172
rect 5165 14112 5229 14116
rect 5245 14172 5309 14176
rect 5245 14116 5249 14172
rect 5249 14116 5305 14172
rect 5305 14116 5309 14172
rect 5245 14112 5309 14116
rect 5325 14172 5389 14176
rect 5325 14116 5329 14172
rect 5329 14116 5385 14172
rect 5385 14116 5389 14172
rect 5325 14112 5389 14116
rect 12031 14172 12095 14176
rect 12031 14116 12035 14172
rect 12035 14116 12091 14172
rect 12091 14116 12095 14172
rect 12031 14112 12095 14116
rect 12111 14172 12175 14176
rect 12111 14116 12115 14172
rect 12115 14116 12171 14172
rect 12171 14116 12175 14172
rect 12111 14112 12175 14116
rect 12191 14172 12255 14176
rect 12191 14116 12195 14172
rect 12195 14116 12251 14172
rect 12251 14116 12255 14172
rect 12191 14112 12255 14116
rect 12271 14172 12335 14176
rect 12271 14116 12275 14172
rect 12275 14116 12331 14172
rect 12331 14116 12335 14172
rect 12271 14112 12335 14116
rect 18977 14172 19041 14176
rect 18977 14116 18981 14172
rect 18981 14116 19037 14172
rect 19037 14116 19041 14172
rect 18977 14112 19041 14116
rect 19057 14172 19121 14176
rect 19057 14116 19061 14172
rect 19061 14116 19117 14172
rect 19117 14116 19121 14172
rect 19057 14112 19121 14116
rect 19137 14172 19201 14176
rect 19137 14116 19141 14172
rect 19141 14116 19197 14172
rect 19197 14116 19201 14172
rect 19137 14112 19201 14116
rect 19217 14172 19281 14176
rect 19217 14116 19221 14172
rect 19221 14116 19277 14172
rect 19277 14116 19281 14172
rect 19217 14112 19281 14116
rect 25923 14172 25987 14176
rect 25923 14116 25927 14172
rect 25927 14116 25983 14172
rect 25983 14116 25987 14172
rect 25923 14112 25987 14116
rect 26003 14172 26067 14176
rect 26003 14116 26007 14172
rect 26007 14116 26063 14172
rect 26063 14116 26067 14172
rect 26003 14112 26067 14116
rect 26083 14172 26147 14176
rect 26083 14116 26087 14172
rect 26087 14116 26143 14172
rect 26143 14116 26147 14172
rect 26083 14112 26147 14116
rect 26163 14172 26227 14176
rect 26163 14116 26167 14172
rect 26167 14116 26223 14172
rect 26223 14116 26227 14172
rect 26163 14112 26227 14116
rect 4425 13628 4489 13632
rect 4425 13572 4429 13628
rect 4429 13572 4485 13628
rect 4485 13572 4489 13628
rect 4425 13568 4489 13572
rect 4505 13628 4569 13632
rect 4505 13572 4509 13628
rect 4509 13572 4565 13628
rect 4565 13572 4569 13628
rect 4505 13568 4569 13572
rect 4585 13628 4649 13632
rect 4585 13572 4589 13628
rect 4589 13572 4645 13628
rect 4645 13572 4649 13628
rect 4585 13568 4649 13572
rect 4665 13628 4729 13632
rect 4665 13572 4669 13628
rect 4669 13572 4725 13628
rect 4725 13572 4729 13628
rect 4665 13568 4729 13572
rect 11371 13628 11435 13632
rect 11371 13572 11375 13628
rect 11375 13572 11431 13628
rect 11431 13572 11435 13628
rect 11371 13568 11435 13572
rect 11451 13628 11515 13632
rect 11451 13572 11455 13628
rect 11455 13572 11511 13628
rect 11511 13572 11515 13628
rect 11451 13568 11515 13572
rect 11531 13628 11595 13632
rect 11531 13572 11535 13628
rect 11535 13572 11591 13628
rect 11591 13572 11595 13628
rect 11531 13568 11595 13572
rect 11611 13628 11675 13632
rect 11611 13572 11615 13628
rect 11615 13572 11671 13628
rect 11671 13572 11675 13628
rect 11611 13568 11675 13572
rect 18317 13628 18381 13632
rect 18317 13572 18321 13628
rect 18321 13572 18377 13628
rect 18377 13572 18381 13628
rect 18317 13568 18381 13572
rect 18397 13628 18461 13632
rect 18397 13572 18401 13628
rect 18401 13572 18457 13628
rect 18457 13572 18461 13628
rect 18397 13568 18461 13572
rect 18477 13628 18541 13632
rect 18477 13572 18481 13628
rect 18481 13572 18537 13628
rect 18537 13572 18541 13628
rect 18477 13568 18541 13572
rect 18557 13628 18621 13632
rect 18557 13572 18561 13628
rect 18561 13572 18617 13628
rect 18617 13572 18621 13628
rect 18557 13568 18621 13572
rect 25263 13628 25327 13632
rect 25263 13572 25267 13628
rect 25267 13572 25323 13628
rect 25323 13572 25327 13628
rect 25263 13568 25327 13572
rect 25343 13628 25407 13632
rect 25343 13572 25347 13628
rect 25347 13572 25403 13628
rect 25403 13572 25407 13628
rect 25343 13568 25407 13572
rect 25423 13628 25487 13632
rect 25423 13572 25427 13628
rect 25427 13572 25483 13628
rect 25483 13572 25487 13628
rect 25423 13568 25487 13572
rect 25503 13628 25567 13632
rect 25503 13572 25507 13628
rect 25507 13572 25563 13628
rect 25563 13572 25567 13628
rect 25503 13568 25567 13572
rect 5085 13084 5149 13088
rect 5085 13028 5089 13084
rect 5089 13028 5145 13084
rect 5145 13028 5149 13084
rect 5085 13024 5149 13028
rect 5165 13084 5229 13088
rect 5165 13028 5169 13084
rect 5169 13028 5225 13084
rect 5225 13028 5229 13084
rect 5165 13024 5229 13028
rect 5245 13084 5309 13088
rect 5245 13028 5249 13084
rect 5249 13028 5305 13084
rect 5305 13028 5309 13084
rect 5245 13024 5309 13028
rect 5325 13084 5389 13088
rect 5325 13028 5329 13084
rect 5329 13028 5385 13084
rect 5385 13028 5389 13084
rect 5325 13024 5389 13028
rect 12031 13084 12095 13088
rect 12031 13028 12035 13084
rect 12035 13028 12091 13084
rect 12091 13028 12095 13084
rect 12031 13024 12095 13028
rect 12111 13084 12175 13088
rect 12111 13028 12115 13084
rect 12115 13028 12171 13084
rect 12171 13028 12175 13084
rect 12111 13024 12175 13028
rect 12191 13084 12255 13088
rect 12191 13028 12195 13084
rect 12195 13028 12251 13084
rect 12251 13028 12255 13084
rect 12191 13024 12255 13028
rect 12271 13084 12335 13088
rect 12271 13028 12275 13084
rect 12275 13028 12331 13084
rect 12331 13028 12335 13084
rect 12271 13024 12335 13028
rect 18977 13084 19041 13088
rect 18977 13028 18981 13084
rect 18981 13028 19037 13084
rect 19037 13028 19041 13084
rect 18977 13024 19041 13028
rect 19057 13084 19121 13088
rect 19057 13028 19061 13084
rect 19061 13028 19117 13084
rect 19117 13028 19121 13084
rect 19057 13024 19121 13028
rect 19137 13084 19201 13088
rect 19137 13028 19141 13084
rect 19141 13028 19197 13084
rect 19197 13028 19201 13084
rect 19137 13024 19201 13028
rect 19217 13084 19281 13088
rect 19217 13028 19221 13084
rect 19221 13028 19277 13084
rect 19277 13028 19281 13084
rect 19217 13024 19281 13028
rect 25923 13084 25987 13088
rect 25923 13028 25927 13084
rect 25927 13028 25983 13084
rect 25983 13028 25987 13084
rect 25923 13024 25987 13028
rect 26003 13084 26067 13088
rect 26003 13028 26007 13084
rect 26007 13028 26063 13084
rect 26063 13028 26067 13084
rect 26003 13024 26067 13028
rect 26083 13084 26147 13088
rect 26083 13028 26087 13084
rect 26087 13028 26143 13084
rect 26143 13028 26147 13084
rect 26083 13024 26147 13028
rect 26163 13084 26227 13088
rect 26163 13028 26167 13084
rect 26167 13028 26223 13084
rect 26223 13028 26227 13084
rect 26163 13024 26227 13028
rect 4425 12540 4489 12544
rect 4425 12484 4429 12540
rect 4429 12484 4485 12540
rect 4485 12484 4489 12540
rect 4425 12480 4489 12484
rect 4505 12540 4569 12544
rect 4505 12484 4509 12540
rect 4509 12484 4565 12540
rect 4565 12484 4569 12540
rect 4505 12480 4569 12484
rect 4585 12540 4649 12544
rect 4585 12484 4589 12540
rect 4589 12484 4645 12540
rect 4645 12484 4649 12540
rect 4585 12480 4649 12484
rect 4665 12540 4729 12544
rect 4665 12484 4669 12540
rect 4669 12484 4725 12540
rect 4725 12484 4729 12540
rect 4665 12480 4729 12484
rect 11371 12540 11435 12544
rect 11371 12484 11375 12540
rect 11375 12484 11431 12540
rect 11431 12484 11435 12540
rect 11371 12480 11435 12484
rect 11451 12540 11515 12544
rect 11451 12484 11455 12540
rect 11455 12484 11511 12540
rect 11511 12484 11515 12540
rect 11451 12480 11515 12484
rect 11531 12540 11595 12544
rect 11531 12484 11535 12540
rect 11535 12484 11591 12540
rect 11591 12484 11595 12540
rect 11531 12480 11595 12484
rect 11611 12540 11675 12544
rect 11611 12484 11615 12540
rect 11615 12484 11671 12540
rect 11671 12484 11675 12540
rect 11611 12480 11675 12484
rect 18317 12540 18381 12544
rect 18317 12484 18321 12540
rect 18321 12484 18377 12540
rect 18377 12484 18381 12540
rect 18317 12480 18381 12484
rect 18397 12540 18461 12544
rect 18397 12484 18401 12540
rect 18401 12484 18457 12540
rect 18457 12484 18461 12540
rect 18397 12480 18461 12484
rect 18477 12540 18541 12544
rect 18477 12484 18481 12540
rect 18481 12484 18537 12540
rect 18537 12484 18541 12540
rect 18477 12480 18541 12484
rect 18557 12540 18621 12544
rect 18557 12484 18561 12540
rect 18561 12484 18617 12540
rect 18617 12484 18621 12540
rect 18557 12480 18621 12484
rect 25263 12540 25327 12544
rect 25263 12484 25267 12540
rect 25267 12484 25323 12540
rect 25323 12484 25327 12540
rect 25263 12480 25327 12484
rect 25343 12540 25407 12544
rect 25343 12484 25347 12540
rect 25347 12484 25403 12540
rect 25403 12484 25407 12540
rect 25343 12480 25407 12484
rect 25423 12540 25487 12544
rect 25423 12484 25427 12540
rect 25427 12484 25483 12540
rect 25483 12484 25487 12540
rect 25423 12480 25487 12484
rect 25503 12540 25567 12544
rect 25503 12484 25507 12540
rect 25507 12484 25563 12540
rect 25563 12484 25567 12540
rect 25503 12480 25567 12484
rect 5085 11996 5149 12000
rect 5085 11940 5089 11996
rect 5089 11940 5145 11996
rect 5145 11940 5149 11996
rect 5085 11936 5149 11940
rect 5165 11996 5229 12000
rect 5165 11940 5169 11996
rect 5169 11940 5225 11996
rect 5225 11940 5229 11996
rect 5165 11936 5229 11940
rect 5245 11996 5309 12000
rect 5245 11940 5249 11996
rect 5249 11940 5305 11996
rect 5305 11940 5309 11996
rect 5245 11936 5309 11940
rect 5325 11996 5389 12000
rect 5325 11940 5329 11996
rect 5329 11940 5385 11996
rect 5385 11940 5389 11996
rect 5325 11936 5389 11940
rect 12031 11996 12095 12000
rect 12031 11940 12035 11996
rect 12035 11940 12091 11996
rect 12091 11940 12095 11996
rect 12031 11936 12095 11940
rect 12111 11996 12175 12000
rect 12111 11940 12115 11996
rect 12115 11940 12171 11996
rect 12171 11940 12175 11996
rect 12111 11936 12175 11940
rect 12191 11996 12255 12000
rect 12191 11940 12195 11996
rect 12195 11940 12251 11996
rect 12251 11940 12255 11996
rect 12191 11936 12255 11940
rect 12271 11996 12335 12000
rect 12271 11940 12275 11996
rect 12275 11940 12331 11996
rect 12331 11940 12335 11996
rect 12271 11936 12335 11940
rect 18977 11996 19041 12000
rect 18977 11940 18981 11996
rect 18981 11940 19037 11996
rect 19037 11940 19041 11996
rect 18977 11936 19041 11940
rect 19057 11996 19121 12000
rect 19057 11940 19061 11996
rect 19061 11940 19117 11996
rect 19117 11940 19121 11996
rect 19057 11936 19121 11940
rect 19137 11996 19201 12000
rect 19137 11940 19141 11996
rect 19141 11940 19197 11996
rect 19197 11940 19201 11996
rect 19137 11936 19201 11940
rect 19217 11996 19281 12000
rect 19217 11940 19221 11996
rect 19221 11940 19277 11996
rect 19277 11940 19281 11996
rect 19217 11936 19281 11940
rect 25923 11996 25987 12000
rect 25923 11940 25927 11996
rect 25927 11940 25983 11996
rect 25983 11940 25987 11996
rect 25923 11936 25987 11940
rect 26003 11996 26067 12000
rect 26003 11940 26007 11996
rect 26007 11940 26063 11996
rect 26063 11940 26067 11996
rect 26003 11936 26067 11940
rect 26083 11996 26147 12000
rect 26083 11940 26087 11996
rect 26087 11940 26143 11996
rect 26143 11940 26147 11996
rect 26083 11936 26147 11940
rect 26163 11996 26227 12000
rect 26163 11940 26167 11996
rect 26167 11940 26223 11996
rect 26223 11940 26227 11996
rect 26163 11936 26227 11940
rect 4425 11452 4489 11456
rect 4425 11396 4429 11452
rect 4429 11396 4485 11452
rect 4485 11396 4489 11452
rect 4425 11392 4489 11396
rect 4505 11452 4569 11456
rect 4505 11396 4509 11452
rect 4509 11396 4565 11452
rect 4565 11396 4569 11452
rect 4505 11392 4569 11396
rect 4585 11452 4649 11456
rect 4585 11396 4589 11452
rect 4589 11396 4645 11452
rect 4645 11396 4649 11452
rect 4585 11392 4649 11396
rect 4665 11452 4729 11456
rect 4665 11396 4669 11452
rect 4669 11396 4725 11452
rect 4725 11396 4729 11452
rect 4665 11392 4729 11396
rect 11371 11452 11435 11456
rect 11371 11396 11375 11452
rect 11375 11396 11431 11452
rect 11431 11396 11435 11452
rect 11371 11392 11435 11396
rect 11451 11452 11515 11456
rect 11451 11396 11455 11452
rect 11455 11396 11511 11452
rect 11511 11396 11515 11452
rect 11451 11392 11515 11396
rect 11531 11452 11595 11456
rect 11531 11396 11535 11452
rect 11535 11396 11591 11452
rect 11591 11396 11595 11452
rect 11531 11392 11595 11396
rect 11611 11452 11675 11456
rect 11611 11396 11615 11452
rect 11615 11396 11671 11452
rect 11671 11396 11675 11452
rect 11611 11392 11675 11396
rect 18317 11452 18381 11456
rect 18317 11396 18321 11452
rect 18321 11396 18377 11452
rect 18377 11396 18381 11452
rect 18317 11392 18381 11396
rect 18397 11452 18461 11456
rect 18397 11396 18401 11452
rect 18401 11396 18457 11452
rect 18457 11396 18461 11452
rect 18397 11392 18461 11396
rect 18477 11452 18541 11456
rect 18477 11396 18481 11452
rect 18481 11396 18537 11452
rect 18537 11396 18541 11452
rect 18477 11392 18541 11396
rect 18557 11452 18621 11456
rect 18557 11396 18561 11452
rect 18561 11396 18617 11452
rect 18617 11396 18621 11452
rect 18557 11392 18621 11396
rect 25263 11452 25327 11456
rect 25263 11396 25267 11452
rect 25267 11396 25323 11452
rect 25323 11396 25327 11452
rect 25263 11392 25327 11396
rect 25343 11452 25407 11456
rect 25343 11396 25347 11452
rect 25347 11396 25403 11452
rect 25403 11396 25407 11452
rect 25343 11392 25407 11396
rect 25423 11452 25487 11456
rect 25423 11396 25427 11452
rect 25427 11396 25483 11452
rect 25483 11396 25487 11452
rect 25423 11392 25487 11396
rect 25503 11452 25567 11456
rect 25503 11396 25507 11452
rect 25507 11396 25563 11452
rect 25563 11396 25567 11452
rect 25503 11392 25567 11396
rect 5085 10908 5149 10912
rect 5085 10852 5089 10908
rect 5089 10852 5145 10908
rect 5145 10852 5149 10908
rect 5085 10848 5149 10852
rect 5165 10908 5229 10912
rect 5165 10852 5169 10908
rect 5169 10852 5225 10908
rect 5225 10852 5229 10908
rect 5165 10848 5229 10852
rect 5245 10908 5309 10912
rect 5245 10852 5249 10908
rect 5249 10852 5305 10908
rect 5305 10852 5309 10908
rect 5245 10848 5309 10852
rect 5325 10908 5389 10912
rect 5325 10852 5329 10908
rect 5329 10852 5385 10908
rect 5385 10852 5389 10908
rect 5325 10848 5389 10852
rect 12031 10908 12095 10912
rect 12031 10852 12035 10908
rect 12035 10852 12091 10908
rect 12091 10852 12095 10908
rect 12031 10848 12095 10852
rect 12111 10908 12175 10912
rect 12111 10852 12115 10908
rect 12115 10852 12171 10908
rect 12171 10852 12175 10908
rect 12111 10848 12175 10852
rect 12191 10908 12255 10912
rect 12191 10852 12195 10908
rect 12195 10852 12251 10908
rect 12251 10852 12255 10908
rect 12191 10848 12255 10852
rect 12271 10908 12335 10912
rect 12271 10852 12275 10908
rect 12275 10852 12331 10908
rect 12331 10852 12335 10908
rect 12271 10848 12335 10852
rect 18977 10908 19041 10912
rect 18977 10852 18981 10908
rect 18981 10852 19037 10908
rect 19037 10852 19041 10908
rect 18977 10848 19041 10852
rect 19057 10908 19121 10912
rect 19057 10852 19061 10908
rect 19061 10852 19117 10908
rect 19117 10852 19121 10908
rect 19057 10848 19121 10852
rect 19137 10908 19201 10912
rect 19137 10852 19141 10908
rect 19141 10852 19197 10908
rect 19197 10852 19201 10908
rect 19137 10848 19201 10852
rect 19217 10908 19281 10912
rect 19217 10852 19221 10908
rect 19221 10852 19277 10908
rect 19277 10852 19281 10908
rect 19217 10848 19281 10852
rect 25923 10908 25987 10912
rect 25923 10852 25927 10908
rect 25927 10852 25983 10908
rect 25983 10852 25987 10908
rect 25923 10848 25987 10852
rect 26003 10908 26067 10912
rect 26003 10852 26007 10908
rect 26007 10852 26063 10908
rect 26063 10852 26067 10908
rect 26003 10848 26067 10852
rect 26083 10908 26147 10912
rect 26083 10852 26087 10908
rect 26087 10852 26143 10908
rect 26143 10852 26147 10908
rect 26083 10848 26147 10852
rect 26163 10908 26227 10912
rect 26163 10852 26167 10908
rect 26167 10852 26223 10908
rect 26223 10852 26227 10908
rect 26163 10848 26227 10852
rect 4425 10364 4489 10368
rect 4425 10308 4429 10364
rect 4429 10308 4485 10364
rect 4485 10308 4489 10364
rect 4425 10304 4489 10308
rect 4505 10364 4569 10368
rect 4505 10308 4509 10364
rect 4509 10308 4565 10364
rect 4565 10308 4569 10364
rect 4505 10304 4569 10308
rect 4585 10364 4649 10368
rect 4585 10308 4589 10364
rect 4589 10308 4645 10364
rect 4645 10308 4649 10364
rect 4585 10304 4649 10308
rect 4665 10364 4729 10368
rect 4665 10308 4669 10364
rect 4669 10308 4725 10364
rect 4725 10308 4729 10364
rect 4665 10304 4729 10308
rect 11371 10364 11435 10368
rect 11371 10308 11375 10364
rect 11375 10308 11431 10364
rect 11431 10308 11435 10364
rect 11371 10304 11435 10308
rect 11451 10364 11515 10368
rect 11451 10308 11455 10364
rect 11455 10308 11511 10364
rect 11511 10308 11515 10364
rect 11451 10304 11515 10308
rect 11531 10364 11595 10368
rect 11531 10308 11535 10364
rect 11535 10308 11591 10364
rect 11591 10308 11595 10364
rect 11531 10304 11595 10308
rect 11611 10364 11675 10368
rect 11611 10308 11615 10364
rect 11615 10308 11671 10364
rect 11671 10308 11675 10364
rect 11611 10304 11675 10308
rect 18317 10364 18381 10368
rect 18317 10308 18321 10364
rect 18321 10308 18377 10364
rect 18377 10308 18381 10364
rect 18317 10304 18381 10308
rect 18397 10364 18461 10368
rect 18397 10308 18401 10364
rect 18401 10308 18457 10364
rect 18457 10308 18461 10364
rect 18397 10304 18461 10308
rect 18477 10364 18541 10368
rect 18477 10308 18481 10364
rect 18481 10308 18537 10364
rect 18537 10308 18541 10364
rect 18477 10304 18541 10308
rect 18557 10364 18621 10368
rect 18557 10308 18561 10364
rect 18561 10308 18617 10364
rect 18617 10308 18621 10364
rect 18557 10304 18621 10308
rect 25263 10364 25327 10368
rect 25263 10308 25267 10364
rect 25267 10308 25323 10364
rect 25323 10308 25327 10364
rect 25263 10304 25327 10308
rect 25343 10364 25407 10368
rect 25343 10308 25347 10364
rect 25347 10308 25403 10364
rect 25403 10308 25407 10364
rect 25343 10304 25407 10308
rect 25423 10364 25487 10368
rect 25423 10308 25427 10364
rect 25427 10308 25483 10364
rect 25483 10308 25487 10364
rect 25423 10304 25487 10308
rect 25503 10364 25567 10368
rect 25503 10308 25507 10364
rect 25507 10308 25563 10364
rect 25563 10308 25567 10364
rect 25503 10304 25567 10308
rect 5085 9820 5149 9824
rect 5085 9764 5089 9820
rect 5089 9764 5145 9820
rect 5145 9764 5149 9820
rect 5085 9760 5149 9764
rect 5165 9820 5229 9824
rect 5165 9764 5169 9820
rect 5169 9764 5225 9820
rect 5225 9764 5229 9820
rect 5165 9760 5229 9764
rect 5245 9820 5309 9824
rect 5245 9764 5249 9820
rect 5249 9764 5305 9820
rect 5305 9764 5309 9820
rect 5245 9760 5309 9764
rect 5325 9820 5389 9824
rect 5325 9764 5329 9820
rect 5329 9764 5385 9820
rect 5385 9764 5389 9820
rect 5325 9760 5389 9764
rect 12031 9820 12095 9824
rect 12031 9764 12035 9820
rect 12035 9764 12091 9820
rect 12091 9764 12095 9820
rect 12031 9760 12095 9764
rect 12111 9820 12175 9824
rect 12111 9764 12115 9820
rect 12115 9764 12171 9820
rect 12171 9764 12175 9820
rect 12111 9760 12175 9764
rect 12191 9820 12255 9824
rect 12191 9764 12195 9820
rect 12195 9764 12251 9820
rect 12251 9764 12255 9820
rect 12191 9760 12255 9764
rect 12271 9820 12335 9824
rect 12271 9764 12275 9820
rect 12275 9764 12331 9820
rect 12331 9764 12335 9820
rect 12271 9760 12335 9764
rect 18977 9820 19041 9824
rect 18977 9764 18981 9820
rect 18981 9764 19037 9820
rect 19037 9764 19041 9820
rect 18977 9760 19041 9764
rect 19057 9820 19121 9824
rect 19057 9764 19061 9820
rect 19061 9764 19117 9820
rect 19117 9764 19121 9820
rect 19057 9760 19121 9764
rect 19137 9820 19201 9824
rect 19137 9764 19141 9820
rect 19141 9764 19197 9820
rect 19197 9764 19201 9820
rect 19137 9760 19201 9764
rect 19217 9820 19281 9824
rect 19217 9764 19221 9820
rect 19221 9764 19277 9820
rect 19277 9764 19281 9820
rect 19217 9760 19281 9764
rect 25923 9820 25987 9824
rect 25923 9764 25927 9820
rect 25927 9764 25983 9820
rect 25983 9764 25987 9820
rect 25923 9760 25987 9764
rect 26003 9820 26067 9824
rect 26003 9764 26007 9820
rect 26007 9764 26063 9820
rect 26063 9764 26067 9820
rect 26003 9760 26067 9764
rect 26083 9820 26147 9824
rect 26083 9764 26087 9820
rect 26087 9764 26143 9820
rect 26143 9764 26147 9820
rect 26083 9760 26147 9764
rect 26163 9820 26227 9824
rect 26163 9764 26167 9820
rect 26167 9764 26223 9820
rect 26223 9764 26227 9820
rect 26163 9760 26227 9764
rect 4425 9276 4489 9280
rect 4425 9220 4429 9276
rect 4429 9220 4485 9276
rect 4485 9220 4489 9276
rect 4425 9216 4489 9220
rect 4505 9276 4569 9280
rect 4505 9220 4509 9276
rect 4509 9220 4565 9276
rect 4565 9220 4569 9276
rect 4505 9216 4569 9220
rect 4585 9276 4649 9280
rect 4585 9220 4589 9276
rect 4589 9220 4645 9276
rect 4645 9220 4649 9276
rect 4585 9216 4649 9220
rect 4665 9276 4729 9280
rect 4665 9220 4669 9276
rect 4669 9220 4725 9276
rect 4725 9220 4729 9276
rect 4665 9216 4729 9220
rect 11371 9276 11435 9280
rect 11371 9220 11375 9276
rect 11375 9220 11431 9276
rect 11431 9220 11435 9276
rect 11371 9216 11435 9220
rect 11451 9276 11515 9280
rect 11451 9220 11455 9276
rect 11455 9220 11511 9276
rect 11511 9220 11515 9276
rect 11451 9216 11515 9220
rect 11531 9276 11595 9280
rect 11531 9220 11535 9276
rect 11535 9220 11591 9276
rect 11591 9220 11595 9276
rect 11531 9216 11595 9220
rect 11611 9276 11675 9280
rect 11611 9220 11615 9276
rect 11615 9220 11671 9276
rect 11671 9220 11675 9276
rect 11611 9216 11675 9220
rect 18317 9276 18381 9280
rect 18317 9220 18321 9276
rect 18321 9220 18377 9276
rect 18377 9220 18381 9276
rect 18317 9216 18381 9220
rect 18397 9276 18461 9280
rect 18397 9220 18401 9276
rect 18401 9220 18457 9276
rect 18457 9220 18461 9276
rect 18397 9216 18461 9220
rect 18477 9276 18541 9280
rect 18477 9220 18481 9276
rect 18481 9220 18537 9276
rect 18537 9220 18541 9276
rect 18477 9216 18541 9220
rect 18557 9276 18621 9280
rect 18557 9220 18561 9276
rect 18561 9220 18617 9276
rect 18617 9220 18621 9276
rect 18557 9216 18621 9220
rect 25263 9276 25327 9280
rect 25263 9220 25267 9276
rect 25267 9220 25323 9276
rect 25323 9220 25327 9276
rect 25263 9216 25327 9220
rect 25343 9276 25407 9280
rect 25343 9220 25347 9276
rect 25347 9220 25403 9276
rect 25403 9220 25407 9276
rect 25343 9216 25407 9220
rect 25423 9276 25487 9280
rect 25423 9220 25427 9276
rect 25427 9220 25483 9276
rect 25483 9220 25487 9276
rect 25423 9216 25487 9220
rect 25503 9276 25567 9280
rect 25503 9220 25507 9276
rect 25507 9220 25563 9276
rect 25563 9220 25567 9276
rect 25503 9216 25567 9220
rect 5085 8732 5149 8736
rect 5085 8676 5089 8732
rect 5089 8676 5145 8732
rect 5145 8676 5149 8732
rect 5085 8672 5149 8676
rect 5165 8732 5229 8736
rect 5165 8676 5169 8732
rect 5169 8676 5225 8732
rect 5225 8676 5229 8732
rect 5165 8672 5229 8676
rect 5245 8732 5309 8736
rect 5245 8676 5249 8732
rect 5249 8676 5305 8732
rect 5305 8676 5309 8732
rect 5245 8672 5309 8676
rect 5325 8732 5389 8736
rect 5325 8676 5329 8732
rect 5329 8676 5385 8732
rect 5385 8676 5389 8732
rect 5325 8672 5389 8676
rect 12031 8732 12095 8736
rect 12031 8676 12035 8732
rect 12035 8676 12091 8732
rect 12091 8676 12095 8732
rect 12031 8672 12095 8676
rect 12111 8732 12175 8736
rect 12111 8676 12115 8732
rect 12115 8676 12171 8732
rect 12171 8676 12175 8732
rect 12111 8672 12175 8676
rect 12191 8732 12255 8736
rect 12191 8676 12195 8732
rect 12195 8676 12251 8732
rect 12251 8676 12255 8732
rect 12191 8672 12255 8676
rect 12271 8732 12335 8736
rect 12271 8676 12275 8732
rect 12275 8676 12331 8732
rect 12331 8676 12335 8732
rect 12271 8672 12335 8676
rect 18977 8732 19041 8736
rect 18977 8676 18981 8732
rect 18981 8676 19037 8732
rect 19037 8676 19041 8732
rect 18977 8672 19041 8676
rect 19057 8732 19121 8736
rect 19057 8676 19061 8732
rect 19061 8676 19117 8732
rect 19117 8676 19121 8732
rect 19057 8672 19121 8676
rect 19137 8732 19201 8736
rect 19137 8676 19141 8732
rect 19141 8676 19197 8732
rect 19197 8676 19201 8732
rect 19137 8672 19201 8676
rect 19217 8732 19281 8736
rect 19217 8676 19221 8732
rect 19221 8676 19277 8732
rect 19277 8676 19281 8732
rect 19217 8672 19281 8676
rect 25923 8732 25987 8736
rect 25923 8676 25927 8732
rect 25927 8676 25983 8732
rect 25983 8676 25987 8732
rect 25923 8672 25987 8676
rect 26003 8732 26067 8736
rect 26003 8676 26007 8732
rect 26007 8676 26063 8732
rect 26063 8676 26067 8732
rect 26003 8672 26067 8676
rect 26083 8732 26147 8736
rect 26083 8676 26087 8732
rect 26087 8676 26143 8732
rect 26143 8676 26147 8732
rect 26083 8672 26147 8676
rect 26163 8732 26227 8736
rect 26163 8676 26167 8732
rect 26167 8676 26223 8732
rect 26223 8676 26227 8732
rect 26163 8672 26227 8676
rect 24900 8196 24964 8260
rect 4425 8188 4489 8192
rect 4425 8132 4429 8188
rect 4429 8132 4485 8188
rect 4485 8132 4489 8188
rect 4425 8128 4489 8132
rect 4505 8188 4569 8192
rect 4505 8132 4509 8188
rect 4509 8132 4565 8188
rect 4565 8132 4569 8188
rect 4505 8128 4569 8132
rect 4585 8188 4649 8192
rect 4585 8132 4589 8188
rect 4589 8132 4645 8188
rect 4645 8132 4649 8188
rect 4585 8128 4649 8132
rect 4665 8188 4729 8192
rect 4665 8132 4669 8188
rect 4669 8132 4725 8188
rect 4725 8132 4729 8188
rect 4665 8128 4729 8132
rect 11371 8188 11435 8192
rect 11371 8132 11375 8188
rect 11375 8132 11431 8188
rect 11431 8132 11435 8188
rect 11371 8128 11435 8132
rect 11451 8188 11515 8192
rect 11451 8132 11455 8188
rect 11455 8132 11511 8188
rect 11511 8132 11515 8188
rect 11451 8128 11515 8132
rect 11531 8188 11595 8192
rect 11531 8132 11535 8188
rect 11535 8132 11591 8188
rect 11591 8132 11595 8188
rect 11531 8128 11595 8132
rect 11611 8188 11675 8192
rect 11611 8132 11615 8188
rect 11615 8132 11671 8188
rect 11671 8132 11675 8188
rect 11611 8128 11675 8132
rect 18317 8188 18381 8192
rect 18317 8132 18321 8188
rect 18321 8132 18377 8188
rect 18377 8132 18381 8188
rect 18317 8128 18381 8132
rect 18397 8188 18461 8192
rect 18397 8132 18401 8188
rect 18401 8132 18457 8188
rect 18457 8132 18461 8188
rect 18397 8128 18461 8132
rect 18477 8188 18541 8192
rect 18477 8132 18481 8188
rect 18481 8132 18537 8188
rect 18537 8132 18541 8188
rect 18477 8128 18541 8132
rect 18557 8188 18621 8192
rect 18557 8132 18561 8188
rect 18561 8132 18617 8188
rect 18617 8132 18621 8188
rect 18557 8128 18621 8132
rect 25263 8188 25327 8192
rect 25263 8132 25267 8188
rect 25267 8132 25323 8188
rect 25323 8132 25327 8188
rect 25263 8128 25327 8132
rect 25343 8188 25407 8192
rect 25343 8132 25347 8188
rect 25347 8132 25403 8188
rect 25403 8132 25407 8188
rect 25343 8128 25407 8132
rect 25423 8188 25487 8192
rect 25423 8132 25427 8188
rect 25427 8132 25483 8188
rect 25483 8132 25487 8188
rect 25423 8128 25487 8132
rect 25503 8188 25567 8192
rect 25503 8132 25507 8188
rect 25507 8132 25563 8188
rect 25563 8132 25567 8188
rect 25503 8128 25567 8132
rect 5085 7644 5149 7648
rect 5085 7588 5089 7644
rect 5089 7588 5145 7644
rect 5145 7588 5149 7644
rect 5085 7584 5149 7588
rect 5165 7644 5229 7648
rect 5165 7588 5169 7644
rect 5169 7588 5225 7644
rect 5225 7588 5229 7644
rect 5165 7584 5229 7588
rect 5245 7644 5309 7648
rect 5245 7588 5249 7644
rect 5249 7588 5305 7644
rect 5305 7588 5309 7644
rect 5245 7584 5309 7588
rect 5325 7644 5389 7648
rect 5325 7588 5329 7644
rect 5329 7588 5385 7644
rect 5385 7588 5389 7644
rect 5325 7584 5389 7588
rect 12031 7644 12095 7648
rect 12031 7588 12035 7644
rect 12035 7588 12091 7644
rect 12091 7588 12095 7644
rect 12031 7584 12095 7588
rect 12111 7644 12175 7648
rect 12111 7588 12115 7644
rect 12115 7588 12171 7644
rect 12171 7588 12175 7644
rect 12111 7584 12175 7588
rect 12191 7644 12255 7648
rect 12191 7588 12195 7644
rect 12195 7588 12251 7644
rect 12251 7588 12255 7644
rect 12191 7584 12255 7588
rect 12271 7644 12335 7648
rect 12271 7588 12275 7644
rect 12275 7588 12331 7644
rect 12331 7588 12335 7644
rect 12271 7584 12335 7588
rect 18977 7644 19041 7648
rect 18977 7588 18981 7644
rect 18981 7588 19037 7644
rect 19037 7588 19041 7644
rect 18977 7584 19041 7588
rect 19057 7644 19121 7648
rect 19057 7588 19061 7644
rect 19061 7588 19117 7644
rect 19117 7588 19121 7644
rect 19057 7584 19121 7588
rect 19137 7644 19201 7648
rect 19137 7588 19141 7644
rect 19141 7588 19197 7644
rect 19197 7588 19201 7644
rect 19137 7584 19201 7588
rect 19217 7644 19281 7648
rect 19217 7588 19221 7644
rect 19221 7588 19277 7644
rect 19277 7588 19281 7644
rect 19217 7584 19281 7588
rect 25923 7644 25987 7648
rect 25923 7588 25927 7644
rect 25927 7588 25983 7644
rect 25983 7588 25987 7644
rect 25923 7584 25987 7588
rect 26003 7644 26067 7648
rect 26003 7588 26007 7644
rect 26007 7588 26063 7644
rect 26063 7588 26067 7644
rect 26003 7584 26067 7588
rect 26083 7644 26147 7648
rect 26083 7588 26087 7644
rect 26087 7588 26143 7644
rect 26143 7588 26147 7644
rect 26083 7584 26147 7588
rect 26163 7644 26227 7648
rect 26163 7588 26167 7644
rect 26167 7588 26223 7644
rect 26223 7588 26227 7644
rect 26163 7584 26227 7588
rect 4425 7100 4489 7104
rect 4425 7044 4429 7100
rect 4429 7044 4485 7100
rect 4485 7044 4489 7100
rect 4425 7040 4489 7044
rect 4505 7100 4569 7104
rect 4505 7044 4509 7100
rect 4509 7044 4565 7100
rect 4565 7044 4569 7100
rect 4505 7040 4569 7044
rect 4585 7100 4649 7104
rect 4585 7044 4589 7100
rect 4589 7044 4645 7100
rect 4645 7044 4649 7100
rect 4585 7040 4649 7044
rect 4665 7100 4729 7104
rect 4665 7044 4669 7100
rect 4669 7044 4725 7100
rect 4725 7044 4729 7100
rect 4665 7040 4729 7044
rect 11371 7100 11435 7104
rect 11371 7044 11375 7100
rect 11375 7044 11431 7100
rect 11431 7044 11435 7100
rect 11371 7040 11435 7044
rect 11451 7100 11515 7104
rect 11451 7044 11455 7100
rect 11455 7044 11511 7100
rect 11511 7044 11515 7100
rect 11451 7040 11515 7044
rect 11531 7100 11595 7104
rect 11531 7044 11535 7100
rect 11535 7044 11591 7100
rect 11591 7044 11595 7100
rect 11531 7040 11595 7044
rect 11611 7100 11675 7104
rect 11611 7044 11615 7100
rect 11615 7044 11671 7100
rect 11671 7044 11675 7100
rect 11611 7040 11675 7044
rect 18317 7100 18381 7104
rect 18317 7044 18321 7100
rect 18321 7044 18377 7100
rect 18377 7044 18381 7100
rect 18317 7040 18381 7044
rect 18397 7100 18461 7104
rect 18397 7044 18401 7100
rect 18401 7044 18457 7100
rect 18457 7044 18461 7100
rect 18397 7040 18461 7044
rect 18477 7100 18541 7104
rect 18477 7044 18481 7100
rect 18481 7044 18537 7100
rect 18537 7044 18541 7100
rect 18477 7040 18541 7044
rect 18557 7100 18621 7104
rect 18557 7044 18561 7100
rect 18561 7044 18617 7100
rect 18617 7044 18621 7100
rect 18557 7040 18621 7044
rect 25263 7100 25327 7104
rect 25263 7044 25267 7100
rect 25267 7044 25323 7100
rect 25323 7044 25327 7100
rect 25263 7040 25327 7044
rect 25343 7100 25407 7104
rect 25343 7044 25347 7100
rect 25347 7044 25403 7100
rect 25403 7044 25407 7100
rect 25343 7040 25407 7044
rect 25423 7100 25487 7104
rect 25423 7044 25427 7100
rect 25427 7044 25483 7100
rect 25483 7044 25487 7100
rect 25423 7040 25487 7044
rect 25503 7100 25567 7104
rect 25503 7044 25507 7100
rect 25507 7044 25563 7100
rect 25563 7044 25567 7100
rect 25503 7040 25567 7044
rect 5085 6556 5149 6560
rect 5085 6500 5089 6556
rect 5089 6500 5145 6556
rect 5145 6500 5149 6556
rect 5085 6496 5149 6500
rect 5165 6556 5229 6560
rect 5165 6500 5169 6556
rect 5169 6500 5225 6556
rect 5225 6500 5229 6556
rect 5165 6496 5229 6500
rect 5245 6556 5309 6560
rect 5245 6500 5249 6556
rect 5249 6500 5305 6556
rect 5305 6500 5309 6556
rect 5245 6496 5309 6500
rect 5325 6556 5389 6560
rect 5325 6500 5329 6556
rect 5329 6500 5385 6556
rect 5385 6500 5389 6556
rect 5325 6496 5389 6500
rect 12031 6556 12095 6560
rect 12031 6500 12035 6556
rect 12035 6500 12091 6556
rect 12091 6500 12095 6556
rect 12031 6496 12095 6500
rect 12111 6556 12175 6560
rect 12111 6500 12115 6556
rect 12115 6500 12171 6556
rect 12171 6500 12175 6556
rect 12111 6496 12175 6500
rect 12191 6556 12255 6560
rect 12191 6500 12195 6556
rect 12195 6500 12251 6556
rect 12251 6500 12255 6556
rect 12191 6496 12255 6500
rect 12271 6556 12335 6560
rect 12271 6500 12275 6556
rect 12275 6500 12331 6556
rect 12331 6500 12335 6556
rect 12271 6496 12335 6500
rect 18977 6556 19041 6560
rect 18977 6500 18981 6556
rect 18981 6500 19037 6556
rect 19037 6500 19041 6556
rect 18977 6496 19041 6500
rect 19057 6556 19121 6560
rect 19057 6500 19061 6556
rect 19061 6500 19117 6556
rect 19117 6500 19121 6556
rect 19057 6496 19121 6500
rect 19137 6556 19201 6560
rect 19137 6500 19141 6556
rect 19141 6500 19197 6556
rect 19197 6500 19201 6556
rect 19137 6496 19201 6500
rect 19217 6556 19281 6560
rect 19217 6500 19221 6556
rect 19221 6500 19277 6556
rect 19277 6500 19281 6556
rect 19217 6496 19281 6500
rect 25923 6556 25987 6560
rect 25923 6500 25927 6556
rect 25927 6500 25983 6556
rect 25983 6500 25987 6556
rect 25923 6496 25987 6500
rect 26003 6556 26067 6560
rect 26003 6500 26007 6556
rect 26007 6500 26063 6556
rect 26063 6500 26067 6556
rect 26003 6496 26067 6500
rect 26083 6556 26147 6560
rect 26083 6500 26087 6556
rect 26087 6500 26143 6556
rect 26143 6500 26147 6556
rect 26083 6496 26147 6500
rect 26163 6556 26227 6560
rect 26163 6500 26167 6556
rect 26167 6500 26223 6556
rect 26223 6500 26227 6556
rect 26163 6496 26227 6500
rect 4425 6012 4489 6016
rect 4425 5956 4429 6012
rect 4429 5956 4485 6012
rect 4485 5956 4489 6012
rect 4425 5952 4489 5956
rect 4505 6012 4569 6016
rect 4505 5956 4509 6012
rect 4509 5956 4565 6012
rect 4565 5956 4569 6012
rect 4505 5952 4569 5956
rect 4585 6012 4649 6016
rect 4585 5956 4589 6012
rect 4589 5956 4645 6012
rect 4645 5956 4649 6012
rect 4585 5952 4649 5956
rect 4665 6012 4729 6016
rect 4665 5956 4669 6012
rect 4669 5956 4725 6012
rect 4725 5956 4729 6012
rect 4665 5952 4729 5956
rect 11371 6012 11435 6016
rect 11371 5956 11375 6012
rect 11375 5956 11431 6012
rect 11431 5956 11435 6012
rect 11371 5952 11435 5956
rect 11451 6012 11515 6016
rect 11451 5956 11455 6012
rect 11455 5956 11511 6012
rect 11511 5956 11515 6012
rect 11451 5952 11515 5956
rect 11531 6012 11595 6016
rect 11531 5956 11535 6012
rect 11535 5956 11591 6012
rect 11591 5956 11595 6012
rect 11531 5952 11595 5956
rect 11611 6012 11675 6016
rect 11611 5956 11615 6012
rect 11615 5956 11671 6012
rect 11671 5956 11675 6012
rect 11611 5952 11675 5956
rect 18317 6012 18381 6016
rect 18317 5956 18321 6012
rect 18321 5956 18377 6012
rect 18377 5956 18381 6012
rect 18317 5952 18381 5956
rect 18397 6012 18461 6016
rect 18397 5956 18401 6012
rect 18401 5956 18457 6012
rect 18457 5956 18461 6012
rect 18397 5952 18461 5956
rect 18477 6012 18541 6016
rect 18477 5956 18481 6012
rect 18481 5956 18537 6012
rect 18537 5956 18541 6012
rect 18477 5952 18541 5956
rect 18557 6012 18621 6016
rect 18557 5956 18561 6012
rect 18561 5956 18617 6012
rect 18617 5956 18621 6012
rect 18557 5952 18621 5956
rect 25263 6012 25327 6016
rect 25263 5956 25267 6012
rect 25267 5956 25323 6012
rect 25323 5956 25327 6012
rect 25263 5952 25327 5956
rect 25343 6012 25407 6016
rect 25343 5956 25347 6012
rect 25347 5956 25403 6012
rect 25403 5956 25407 6012
rect 25343 5952 25407 5956
rect 25423 6012 25487 6016
rect 25423 5956 25427 6012
rect 25427 5956 25483 6012
rect 25483 5956 25487 6012
rect 25423 5952 25487 5956
rect 25503 6012 25567 6016
rect 25503 5956 25507 6012
rect 25507 5956 25563 6012
rect 25563 5956 25567 6012
rect 25503 5952 25567 5956
rect 5085 5468 5149 5472
rect 5085 5412 5089 5468
rect 5089 5412 5145 5468
rect 5145 5412 5149 5468
rect 5085 5408 5149 5412
rect 5165 5468 5229 5472
rect 5165 5412 5169 5468
rect 5169 5412 5225 5468
rect 5225 5412 5229 5468
rect 5165 5408 5229 5412
rect 5245 5468 5309 5472
rect 5245 5412 5249 5468
rect 5249 5412 5305 5468
rect 5305 5412 5309 5468
rect 5245 5408 5309 5412
rect 5325 5468 5389 5472
rect 5325 5412 5329 5468
rect 5329 5412 5385 5468
rect 5385 5412 5389 5468
rect 5325 5408 5389 5412
rect 12031 5468 12095 5472
rect 12031 5412 12035 5468
rect 12035 5412 12091 5468
rect 12091 5412 12095 5468
rect 12031 5408 12095 5412
rect 12111 5468 12175 5472
rect 12111 5412 12115 5468
rect 12115 5412 12171 5468
rect 12171 5412 12175 5468
rect 12111 5408 12175 5412
rect 12191 5468 12255 5472
rect 12191 5412 12195 5468
rect 12195 5412 12251 5468
rect 12251 5412 12255 5468
rect 12191 5408 12255 5412
rect 12271 5468 12335 5472
rect 12271 5412 12275 5468
rect 12275 5412 12331 5468
rect 12331 5412 12335 5468
rect 12271 5408 12335 5412
rect 18977 5468 19041 5472
rect 18977 5412 18981 5468
rect 18981 5412 19037 5468
rect 19037 5412 19041 5468
rect 18977 5408 19041 5412
rect 19057 5468 19121 5472
rect 19057 5412 19061 5468
rect 19061 5412 19117 5468
rect 19117 5412 19121 5468
rect 19057 5408 19121 5412
rect 19137 5468 19201 5472
rect 19137 5412 19141 5468
rect 19141 5412 19197 5468
rect 19197 5412 19201 5468
rect 19137 5408 19201 5412
rect 19217 5468 19281 5472
rect 19217 5412 19221 5468
rect 19221 5412 19277 5468
rect 19277 5412 19281 5468
rect 19217 5408 19281 5412
rect 25923 5468 25987 5472
rect 25923 5412 25927 5468
rect 25927 5412 25983 5468
rect 25983 5412 25987 5468
rect 25923 5408 25987 5412
rect 26003 5468 26067 5472
rect 26003 5412 26007 5468
rect 26007 5412 26063 5468
rect 26063 5412 26067 5468
rect 26003 5408 26067 5412
rect 26083 5468 26147 5472
rect 26083 5412 26087 5468
rect 26087 5412 26143 5468
rect 26143 5412 26147 5468
rect 26083 5408 26147 5412
rect 26163 5468 26227 5472
rect 26163 5412 26167 5468
rect 26167 5412 26223 5468
rect 26223 5412 26227 5468
rect 26163 5408 26227 5412
rect 4425 4924 4489 4928
rect 4425 4868 4429 4924
rect 4429 4868 4485 4924
rect 4485 4868 4489 4924
rect 4425 4864 4489 4868
rect 4505 4924 4569 4928
rect 4505 4868 4509 4924
rect 4509 4868 4565 4924
rect 4565 4868 4569 4924
rect 4505 4864 4569 4868
rect 4585 4924 4649 4928
rect 4585 4868 4589 4924
rect 4589 4868 4645 4924
rect 4645 4868 4649 4924
rect 4585 4864 4649 4868
rect 4665 4924 4729 4928
rect 4665 4868 4669 4924
rect 4669 4868 4725 4924
rect 4725 4868 4729 4924
rect 4665 4864 4729 4868
rect 11371 4924 11435 4928
rect 11371 4868 11375 4924
rect 11375 4868 11431 4924
rect 11431 4868 11435 4924
rect 11371 4864 11435 4868
rect 11451 4924 11515 4928
rect 11451 4868 11455 4924
rect 11455 4868 11511 4924
rect 11511 4868 11515 4924
rect 11451 4864 11515 4868
rect 11531 4924 11595 4928
rect 11531 4868 11535 4924
rect 11535 4868 11591 4924
rect 11591 4868 11595 4924
rect 11531 4864 11595 4868
rect 11611 4924 11675 4928
rect 11611 4868 11615 4924
rect 11615 4868 11671 4924
rect 11671 4868 11675 4924
rect 11611 4864 11675 4868
rect 18317 4924 18381 4928
rect 18317 4868 18321 4924
rect 18321 4868 18377 4924
rect 18377 4868 18381 4924
rect 18317 4864 18381 4868
rect 18397 4924 18461 4928
rect 18397 4868 18401 4924
rect 18401 4868 18457 4924
rect 18457 4868 18461 4924
rect 18397 4864 18461 4868
rect 18477 4924 18541 4928
rect 18477 4868 18481 4924
rect 18481 4868 18537 4924
rect 18537 4868 18541 4924
rect 18477 4864 18541 4868
rect 18557 4924 18621 4928
rect 18557 4868 18561 4924
rect 18561 4868 18617 4924
rect 18617 4868 18621 4924
rect 18557 4864 18621 4868
rect 25263 4924 25327 4928
rect 25263 4868 25267 4924
rect 25267 4868 25323 4924
rect 25323 4868 25327 4924
rect 25263 4864 25327 4868
rect 25343 4924 25407 4928
rect 25343 4868 25347 4924
rect 25347 4868 25403 4924
rect 25403 4868 25407 4924
rect 25343 4864 25407 4868
rect 25423 4924 25487 4928
rect 25423 4868 25427 4924
rect 25427 4868 25483 4924
rect 25483 4868 25487 4924
rect 25423 4864 25487 4868
rect 25503 4924 25567 4928
rect 25503 4868 25507 4924
rect 25507 4868 25563 4924
rect 25563 4868 25567 4924
rect 25503 4864 25567 4868
rect 5085 4380 5149 4384
rect 5085 4324 5089 4380
rect 5089 4324 5145 4380
rect 5145 4324 5149 4380
rect 5085 4320 5149 4324
rect 5165 4380 5229 4384
rect 5165 4324 5169 4380
rect 5169 4324 5225 4380
rect 5225 4324 5229 4380
rect 5165 4320 5229 4324
rect 5245 4380 5309 4384
rect 5245 4324 5249 4380
rect 5249 4324 5305 4380
rect 5305 4324 5309 4380
rect 5245 4320 5309 4324
rect 5325 4380 5389 4384
rect 5325 4324 5329 4380
rect 5329 4324 5385 4380
rect 5385 4324 5389 4380
rect 5325 4320 5389 4324
rect 12031 4380 12095 4384
rect 12031 4324 12035 4380
rect 12035 4324 12091 4380
rect 12091 4324 12095 4380
rect 12031 4320 12095 4324
rect 12111 4380 12175 4384
rect 12111 4324 12115 4380
rect 12115 4324 12171 4380
rect 12171 4324 12175 4380
rect 12111 4320 12175 4324
rect 12191 4380 12255 4384
rect 12191 4324 12195 4380
rect 12195 4324 12251 4380
rect 12251 4324 12255 4380
rect 12191 4320 12255 4324
rect 12271 4380 12335 4384
rect 12271 4324 12275 4380
rect 12275 4324 12331 4380
rect 12331 4324 12335 4380
rect 12271 4320 12335 4324
rect 18977 4380 19041 4384
rect 18977 4324 18981 4380
rect 18981 4324 19037 4380
rect 19037 4324 19041 4380
rect 18977 4320 19041 4324
rect 19057 4380 19121 4384
rect 19057 4324 19061 4380
rect 19061 4324 19117 4380
rect 19117 4324 19121 4380
rect 19057 4320 19121 4324
rect 19137 4380 19201 4384
rect 19137 4324 19141 4380
rect 19141 4324 19197 4380
rect 19197 4324 19201 4380
rect 19137 4320 19201 4324
rect 19217 4380 19281 4384
rect 19217 4324 19221 4380
rect 19221 4324 19277 4380
rect 19277 4324 19281 4380
rect 19217 4320 19281 4324
rect 25923 4380 25987 4384
rect 25923 4324 25927 4380
rect 25927 4324 25983 4380
rect 25983 4324 25987 4380
rect 25923 4320 25987 4324
rect 26003 4380 26067 4384
rect 26003 4324 26007 4380
rect 26007 4324 26063 4380
rect 26063 4324 26067 4380
rect 26003 4320 26067 4324
rect 26083 4380 26147 4384
rect 26083 4324 26087 4380
rect 26087 4324 26143 4380
rect 26143 4324 26147 4380
rect 26083 4320 26147 4324
rect 26163 4380 26227 4384
rect 26163 4324 26167 4380
rect 26167 4324 26223 4380
rect 26223 4324 26227 4380
rect 26163 4320 26227 4324
rect 4425 3836 4489 3840
rect 4425 3780 4429 3836
rect 4429 3780 4485 3836
rect 4485 3780 4489 3836
rect 4425 3776 4489 3780
rect 4505 3836 4569 3840
rect 4505 3780 4509 3836
rect 4509 3780 4565 3836
rect 4565 3780 4569 3836
rect 4505 3776 4569 3780
rect 4585 3836 4649 3840
rect 4585 3780 4589 3836
rect 4589 3780 4645 3836
rect 4645 3780 4649 3836
rect 4585 3776 4649 3780
rect 4665 3836 4729 3840
rect 4665 3780 4669 3836
rect 4669 3780 4725 3836
rect 4725 3780 4729 3836
rect 4665 3776 4729 3780
rect 11371 3836 11435 3840
rect 11371 3780 11375 3836
rect 11375 3780 11431 3836
rect 11431 3780 11435 3836
rect 11371 3776 11435 3780
rect 11451 3836 11515 3840
rect 11451 3780 11455 3836
rect 11455 3780 11511 3836
rect 11511 3780 11515 3836
rect 11451 3776 11515 3780
rect 11531 3836 11595 3840
rect 11531 3780 11535 3836
rect 11535 3780 11591 3836
rect 11591 3780 11595 3836
rect 11531 3776 11595 3780
rect 11611 3836 11675 3840
rect 11611 3780 11615 3836
rect 11615 3780 11671 3836
rect 11671 3780 11675 3836
rect 11611 3776 11675 3780
rect 18317 3836 18381 3840
rect 18317 3780 18321 3836
rect 18321 3780 18377 3836
rect 18377 3780 18381 3836
rect 18317 3776 18381 3780
rect 18397 3836 18461 3840
rect 18397 3780 18401 3836
rect 18401 3780 18457 3836
rect 18457 3780 18461 3836
rect 18397 3776 18461 3780
rect 18477 3836 18541 3840
rect 18477 3780 18481 3836
rect 18481 3780 18537 3836
rect 18537 3780 18541 3836
rect 18477 3776 18541 3780
rect 18557 3836 18621 3840
rect 18557 3780 18561 3836
rect 18561 3780 18617 3836
rect 18617 3780 18621 3836
rect 18557 3776 18621 3780
rect 25263 3836 25327 3840
rect 25263 3780 25267 3836
rect 25267 3780 25323 3836
rect 25323 3780 25327 3836
rect 25263 3776 25327 3780
rect 25343 3836 25407 3840
rect 25343 3780 25347 3836
rect 25347 3780 25403 3836
rect 25403 3780 25407 3836
rect 25343 3776 25407 3780
rect 25423 3836 25487 3840
rect 25423 3780 25427 3836
rect 25427 3780 25483 3836
rect 25483 3780 25487 3836
rect 25423 3776 25487 3780
rect 25503 3836 25567 3840
rect 25503 3780 25507 3836
rect 25507 3780 25563 3836
rect 25563 3780 25567 3836
rect 25503 3776 25567 3780
rect 5085 3292 5149 3296
rect 5085 3236 5089 3292
rect 5089 3236 5145 3292
rect 5145 3236 5149 3292
rect 5085 3232 5149 3236
rect 5165 3292 5229 3296
rect 5165 3236 5169 3292
rect 5169 3236 5225 3292
rect 5225 3236 5229 3292
rect 5165 3232 5229 3236
rect 5245 3292 5309 3296
rect 5245 3236 5249 3292
rect 5249 3236 5305 3292
rect 5305 3236 5309 3292
rect 5245 3232 5309 3236
rect 5325 3292 5389 3296
rect 5325 3236 5329 3292
rect 5329 3236 5385 3292
rect 5385 3236 5389 3292
rect 5325 3232 5389 3236
rect 12031 3292 12095 3296
rect 12031 3236 12035 3292
rect 12035 3236 12091 3292
rect 12091 3236 12095 3292
rect 12031 3232 12095 3236
rect 12111 3292 12175 3296
rect 12111 3236 12115 3292
rect 12115 3236 12171 3292
rect 12171 3236 12175 3292
rect 12111 3232 12175 3236
rect 12191 3292 12255 3296
rect 12191 3236 12195 3292
rect 12195 3236 12251 3292
rect 12251 3236 12255 3292
rect 12191 3232 12255 3236
rect 12271 3292 12335 3296
rect 12271 3236 12275 3292
rect 12275 3236 12331 3292
rect 12331 3236 12335 3292
rect 12271 3232 12335 3236
rect 18977 3292 19041 3296
rect 18977 3236 18981 3292
rect 18981 3236 19037 3292
rect 19037 3236 19041 3292
rect 18977 3232 19041 3236
rect 19057 3292 19121 3296
rect 19057 3236 19061 3292
rect 19061 3236 19117 3292
rect 19117 3236 19121 3292
rect 19057 3232 19121 3236
rect 19137 3292 19201 3296
rect 19137 3236 19141 3292
rect 19141 3236 19197 3292
rect 19197 3236 19201 3292
rect 19137 3232 19201 3236
rect 19217 3292 19281 3296
rect 19217 3236 19221 3292
rect 19221 3236 19277 3292
rect 19277 3236 19281 3292
rect 19217 3232 19281 3236
rect 25923 3292 25987 3296
rect 25923 3236 25927 3292
rect 25927 3236 25983 3292
rect 25983 3236 25987 3292
rect 25923 3232 25987 3236
rect 26003 3292 26067 3296
rect 26003 3236 26007 3292
rect 26007 3236 26063 3292
rect 26063 3236 26067 3292
rect 26003 3232 26067 3236
rect 26083 3292 26147 3296
rect 26083 3236 26087 3292
rect 26087 3236 26143 3292
rect 26143 3236 26147 3292
rect 26083 3232 26147 3236
rect 26163 3292 26227 3296
rect 26163 3236 26167 3292
rect 26167 3236 26223 3292
rect 26223 3236 26227 3292
rect 26163 3232 26227 3236
rect 4425 2748 4489 2752
rect 4425 2692 4429 2748
rect 4429 2692 4485 2748
rect 4485 2692 4489 2748
rect 4425 2688 4489 2692
rect 4505 2748 4569 2752
rect 4505 2692 4509 2748
rect 4509 2692 4565 2748
rect 4565 2692 4569 2748
rect 4505 2688 4569 2692
rect 4585 2748 4649 2752
rect 4585 2692 4589 2748
rect 4589 2692 4645 2748
rect 4645 2692 4649 2748
rect 4585 2688 4649 2692
rect 4665 2748 4729 2752
rect 4665 2692 4669 2748
rect 4669 2692 4725 2748
rect 4725 2692 4729 2748
rect 4665 2688 4729 2692
rect 11371 2748 11435 2752
rect 11371 2692 11375 2748
rect 11375 2692 11431 2748
rect 11431 2692 11435 2748
rect 11371 2688 11435 2692
rect 11451 2748 11515 2752
rect 11451 2692 11455 2748
rect 11455 2692 11511 2748
rect 11511 2692 11515 2748
rect 11451 2688 11515 2692
rect 11531 2748 11595 2752
rect 11531 2692 11535 2748
rect 11535 2692 11591 2748
rect 11591 2692 11595 2748
rect 11531 2688 11595 2692
rect 11611 2748 11675 2752
rect 11611 2692 11615 2748
rect 11615 2692 11671 2748
rect 11671 2692 11675 2748
rect 11611 2688 11675 2692
rect 18317 2748 18381 2752
rect 18317 2692 18321 2748
rect 18321 2692 18377 2748
rect 18377 2692 18381 2748
rect 18317 2688 18381 2692
rect 18397 2748 18461 2752
rect 18397 2692 18401 2748
rect 18401 2692 18457 2748
rect 18457 2692 18461 2748
rect 18397 2688 18461 2692
rect 18477 2748 18541 2752
rect 18477 2692 18481 2748
rect 18481 2692 18537 2748
rect 18537 2692 18541 2748
rect 18477 2688 18541 2692
rect 18557 2748 18621 2752
rect 18557 2692 18561 2748
rect 18561 2692 18617 2748
rect 18617 2692 18621 2748
rect 18557 2688 18621 2692
rect 25263 2748 25327 2752
rect 25263 2692 25267 2748
rect 25267 2692 25323 2748
rect 25323 2692 25327 2748
rect 25263 2688 25327 2692
rect 25343 2748 25407 2752
rect 25343 2692 25347 2748
rect 25347 2692 25403 2748
rect 25403 2692 25407 2748
rect 25343 2688 25407 2692
rect 25423 2748 25487 2752
rect 25423 2692 25427 2748
rect 25427 2692 25483 2748
rect 25483 2692 25487 2748
rect 25423 2688 25487 2692
rect 25503 2748 25567 2752
rect 25503 2692 25507 2748
rect 25507 2692 25563 2748
rect 25563 2692 25567 2748
rect 25503 2688 25567 2692
rect 5085 2204 5149 2208
rect 5085 2148 5089 2204
rect 5089 2148 5145 2204
rect 5145 2148 5149 2204
rect 5085 2144 5149 2148
rect 5165 2204 5229 2208
rect 5165 2148 5169 2204
rect 5169 2148 5225 2204
rect 5225 2148 5229 2204
rect 5165 2144 5229 2148
rect 5245 2204 5309 2208
rect 5245 2148 5249 2204
rect 5249 2148 5305 2204
rect 5305 2148 5309 2204
rect 5245 2144 5309 2148
rect 5325 2204 5389 2208
rect 5325 2148 5329 2204
rect 5329 2148 5385 2204
rect 5385 2148 5389 2204
rect 5325 2144 5389 2148
rect 12031 2204 12095 2208
rect 12031 2148 12035 2204
rect 12035 2148 12091 2204
rect 12091 2148 12095 2204
rect 12031 2144 12095 2148
rect 12111 2204 12175 2208
rect 12111 2148 12115 2204
rect 12115 2148 12171 2204
rect 12171 2148 12175 2204
rect 12111 2144 12175 2148
rect 12191 2204 12255 2208
rect 12191 2148 12195 2204
rect 12195 2148 12251 2204
rect 12251 2148 12255 2204
rect 12191 2144 12255 2148
rect 12271 2204 12335 2208
rect 12271 2148 12275 2204
rect 12275 2148 12331 2204
rect 12331 2148 12335 2204
rect 12271 2144 12335 2148
rect 18977 2204 19041 2208
rect 18977 2148 18981 2204
rect 18981 2148 19037 2204
rect 19037 2148 19041 2204
rect 18977 2144 19041 2148
rect 19057 2204 19121 2208
rect 19057 2148 19061 2204
rect 19061 2148 19117 2204
rect 19117 2148 19121 2204
rect 19057 2144 19121 2148
rect 19137 2204 19201 2208
rect 19137 2148 19141 2204
rect 19141 2148 19197 2204
rect 19197 2148 19201 2204
rect 19137 2144 19201 2148
rect 19217 2204 19281 2208
rect 19217 2148 19221 2204
rect 19221 2148 19277 2204
rect 19277 2148 19281 2204
rect 19217 2144 19281 2148
rect 25923 2204 25987 2208
rect 25923 2148 25927 2204
rect 25927 2148 25983 2204
rect 25983 2148 25987 2204
rect 25923 2144 25987 2148
rect 26003 2204 26067 2208
rect 26003 2148 26007 2204
rect 26007 2148 26063 2204
rect 26063 2148 26067 2204
rect 26003 2144 26067 2148
rect 26083 2204 26147 2208
rect 26083 2148 26087 2204
rect 26087 2148 26143 2204
rect 26143 2148 26147 2204
rect 26083 2144 26147 2148
rect 26163 2204 26227 2208
rect 26163 2148 26167 2204
rect 26167 2148 26223 2204
rect 26223 2148 26227 2204
rect 26163 2144 26227 2148
<< metal4 >>
rect 4417 27776 4737 27792
rect 4417 27712 4425 27776
rect 4489 27712 4505 27776
rect 4569 27712 4585 27776
rect 4649 27712 4665 27776
rect 4729 27712 4737 27776
rect 4417 26688 4737 27712
rect 4417 26624 4425 26688
rect 4489 26624 4505 26688
rect 4569 26624 4585 26688
rect 4649 26624 4665 26688
rect 4729 26624 4737 26688
rect 4417 25600 4737 26624
rect 4417 25536 4425 25600
rect 4489 25536 4505 25600
rect 4569 25536 4585 25600
rect 4649 25536 4665 25600
rect 4729 25536 4737 25600
rect 4417 24666 4737 25536
rect 4417 24512 4459 24666
rect 4695 24512 4737 24666
rect 4417 24448 4425 24512
rect 4729 24448 4737 24512
rect 4417 24430 4459 24448
rect 4695 24430 4737 24448
rect 4417 23424 4737 24430
rect 4417 23360 4425 23424
rect 4489 23360 4505 23424
rect 4569 23360 4585 23424
rect 4649 23360 4665 23424
rect 4729 23360 4737 23424
rect 4417 22336 4737 23360
rect 4417 22272 4425 22336
rect 4489 22272 4505 22336
rect 4569 22272 4585 22336
rect 4649 22272 4665 22336
rect 4729 22272 4737 22336
rect 4417 21248 4737 22272
rect 4417 21184 4425 21248
rect 4489 21184 4505 21248
rect 4569 21184 4585 21248
rect 4649 21184 4665 21248
rect 4729 21184 4737 21248
rect 4417 20160 4737 21184
rect 4417 20096 4425 20160
rect 4489 20096 4505 20160
rect 4569 20096 4585 20160
rect 4649 20096 4665 20160
rect 4729 20096 4737 20160
rect 4417 19072 4737 20096
rect 4417 19008 4425 19072
rect 4489 19008 4505 19072
rect 4569 19008 4585 19072
rect 4649 19008 4665 19072
rect 4729 19008 4737 19072
rect 4417 18274 4737 19008
rect 4417 18038 4459 18274
rect 4695 18038 4737 18274
rect 4417 17984 4737 18038
rect 4417 17920 4425 17984
rect 4489 17920 4505 17984
rect 4569 17920 4585 17984
rect 4649 17920 4665 17984
rect 4729 17920 4737 17984
rect 4417 16896 4737 17920
rect 4417 16832 4425 16896
rect 4489 16832 4505 16896
rect 4569 16832 4585 16896
rect 4649 16832 4665 16896
rect 4729 16832 4737 16896
rect 4417 15808 4737 16832
rect 4417 15744 4425 15808
rect 4489 15744 4505 15808
rect 4569 15744 4585 15808
rect 4649 15744 4665 15808
rect 4729 15744 4737 15808
rect 4417 14720 4737 15744
rect 4417 14656 4425 14720
rect 4489 14656 4505 14720
rect 4569 14656 4585 14720
rect 4649 14656 4665 14720
rect 4729 14656 4737 14720
rect 4417 13632 4737 14656
rect 4417 13568 4425 13632
rect 4489 13568 4505 13632
rect 4569 13568 4585 13632
rect 4649 13568 4665 13632
rect 4729 13568 4737 13632
rect 4417 12544 4737 13568
rect 4417 12480 4425 12544
rect 4489 12480 4505 12544
rect 4569 12480 4585 12544
rect 4649 12480 4665 12544
rect 4729 12480 4737 12544
rect 4417 11882 4737 12480
rect 4417 11646 4459 11882
rect 4695 11646 4737 11882
rect 4417 11456 4737 11646
rect 4417 11392 4425 11456
rect 4489 11392 4505 11456
rect 4569 11392 4585 11456
rect 4649 11392 4665 11456
rect 4729 11392 4737 11456
rect 4417 10368 4737 11392
rect 4417 10304 4425 10368
rect 4489 10304 4505 10368
rect 4569 10304 4585 10368
rect 4649 10304 4665 10368
rect 4729 10304 4737 10368
rect 4417 9280 4737 10304
rect 4417 9216 4425 9280
rect 4489 9216 4505 9280
rect 4569 9216 4585 9280
rect 4649 9216 4665 9280
rect 4729 9216 4737 9280
rect 4417 8192 4737 9216
rect 4417 8128 4425 8192
rect 4489 8128 4505 8192
rect 4569 8128 4585 8192
rect 4649 8128 4665 8192
rect 4729 8128 4737 8192
rect 4417 7104 4737 8128
rect 4417 7040 4425 7104
rect 4489 7040 4505 7104
rect 4569 7040 4585 7104
rect 4649 7040 4665 7104
rect 4729 7040 4737 7104
rect 4417 6016 4737 7040
rect 4417 5952 4425 6016
rect 4489 5952 4505 6016
rect 4569 5952 4585 6016
rect 4649 5952 4665 6016
rect 4729 5952 4737 6016
rect 4417 5490 4737 5952
rect 4417 5254 4459 5490
rect 4695 5254 4737 5490
rect 4417 4928 4737 5254
rect 4417 4864 4425 4928
rect 4489 4864 4505 4928
rect 4569 4864 4585 4928
rect 4649 4864 4665 4928
rect 4729 4864 4737 4928
rect 4417 3840 4737 4864
rect 4417 3776 4425 3840
rect 4489 3776 4505 3840
rect 4569 3776 4585 3840
rect 4649 3776 4665 3840
rect 4729 3776 4737 3840
rect 4417 2752 4737 3776
rect 4417 2688 4425 2752
rect 4489 2688 4505 2752
rect 4569 2688 4585 2752
rect 4649 2688 4665 2752
rect 4729 2688 4737 2752
rect 4417 2128 4737 2688
rect 5077 27232 5397 27792
rect 5077 27168 5085 27232
rect 5149 27168 5165 27232
rect 5229 27168 5245 27232
rect 5309 27168 5325 27232
rect 5389 27168 5397 27232
rect 5077 26144 5397 27168
rect 5077 26080 5085 26144
rect 5149 26080 5165 26144
rect 5229 26080 5245 26144
rect 5309 26080 5325 26144
rect 5389 26080 5397 26144
rect 5077 25326 5397 26080
rect 5077 25090 5119 25326
rect 5355 25090 5397 25326
rect 5077 25056 5397 25090
rect 5077 24992 5085 25056
rect 5149 24992 5165 25056
rect 5229 24992 5245 25056
rect 5309 24992 5325 25056
rect 5389 24992 5397 25056
rect 5077 23968 5397 24992
rect 5077 23904 5085 23968
rect 5149 23904 5165 23968
rect 5229 23904 5245 23968
rect 5309 23904 5325 23968
rect 5389 23904 5397 23968
rect 5077 22880 5397 23904
rect 5077 22816 5085 22880
rect 5149 22816 5165 22880
rect 5229 22816 5245 22880
rect 5309 22816 5325 22880
rect 5389 22816 5397 22880
rect 5077 21792 5397 22816
rect 5077 21728 5085 21792
rect 5149 21728 5165 21792
rect 5229 21728 5245 21792
rect 5309 21728 5325 21792
rect 5389 21728 5397 21792
rect 5077 20704 5397 21728
rect 5077 20640 5085 20704
rect 5149 20640 5165 20704
rect 5229 20640 5245 20704
rect 5309 20640 5325 20704
rect 5389 20640 5397 20704
rect 5077 19616 5397 20640
rect 5077 19552 5085 19616
rect 5149 19552 5165 19616
rect 5229 19552 5245 19616
rect 5309 19552 5325 19616
rect 5389 19552 5397 19616
rect 5077 18934 5397 19552
rect 5077 18698 5119 18934
rect 5355 18698 5397 18934
rect 5077 18528 5397 18698
rect 5077 18464 5085 18528
rect 5149 18464 5165 18528
rect 5229 18464 5245 18528
rect 5309 18464 5325 18528
rect 5389 18464 5397 18528
rect 5077 17440 5397 18464
rect 5077 17376 5085 17440
rect 5149 17376 5165 17440
rect 5229 17376 5245 17440
rect 5309 17376 5325 17440
rect 5389 17376 5397 17440
rect 5077 16352 5397 17376
rect 5077 16288 5085 16352
rect 5149 16288 5165 16352
rect 5229 16288 5245 16352
rect 5309 16288 5325 16352
rect 5389 16288 5397 16352
rect 5077 15264 5397 16288
rect 5077 15200 5085 15264
rect 5149 15200 5165 15264
rect 5229 15200 5245 15264
rect 5309 15200 5325 15264
rect 5389 15200 5397 15264
rect 5077 14176 5397 15200
rect 5077 14112 5085 14176
rect 5149 14112 5165 14176
rect 5229 14112 5245 14176
rect 5309 14112 5325 14176
rect 5389 14112 5397 14176
rect 5077 13088 5397 14112
rect 5077 13024 5085 13088
rect 5149 13024 5165 13088
rect 5229 13024 5245 13088
rect 5309 13024 5325 13088
rect 5389 13024 5397 13088
rect 5077 12542 5397 13024
rect 5077 12306 5119 12542
rect 5355 12306 5397 12542
rect 5077 12000 5397 12306
rect 5077 11936 5085 12000
rect 5149 11936 5165 12000
rect 5229 11936 5245 12000
rect 5309 11936 5325 12000
rect 5389 11936 5397 12000
rect 5077 10912 5397 11936
rect 5077 10848 5085 10912
rect 5149 10848 5165 10912
rect 5229 10848 5245 10912
rect 5309 10848 5325 10912
rect 5389 10848 5397 10912
rect 5077 9824 5397 10848
rect 5077 9760 5085 9824
rect 5149 9760 5165 9824
rect 5229 9760 5245 9824
rect 5309 9760 5325 9824
rect 5389 9760 5397 9824
rect 5077 8736 5397 9760
rect 5077 8672 5085 8736
rect 5149 8672 5165 8736
rect 5229 8672 5245 8736
rect 5309 8672 5325 8736
rect 5389 8672 5397 8736
rect 5077 7648 5397 8672
rect 5077 7584 5085 7648
rect 5149 7584 5165 7648
rect 5229 7584 5245 7648
rect 5309 7584 5325 7648
rect 5389 7584 5397 7648
rect 5077 6560 5397 7584
rect 5077 6496 5085 6560
rect 5149 6496 5165 6560
rect 5229 6496 5245 6560
rect 5309 6496 5325 6560
rect 5389 6496 5397 6560
rect 5077 6150 5397 6496
rect 5077 5914 5119 6150
rect 5355 5914 5397 6150
rect 5077 5472 5397 5914
rect 5077 5408 5085 5472
rect 5149 5408 5165 5472
rect 5229 5408 5245 5472
rect 5309 5408 5325 5472
rect 5389 5408 5397 5472
rect 5077 4384 5397 5408
rect 5077 4320 5085 4384
rect 5149 4320 5165 4384
rect 5229 4320 5245 4384
rect 5309 4320 5325 4384
rect 5389 4320 5397 4384
rect 5077 3296 5397 4320
rect 5077 3232 5085 3296
rect 5149 3232 5165 3296
rect 5229 3232 5245 3296
rect 5309 3232 5325 3296
rect 5389 3232 5397 3296
rect 5077 2208 5397 3232
rect 5077 2144 5085 2208
rect 5149 2144 5165 2208
rect 5229 2144 5245 2208
rect 5309 2144 5325 2208
rect 5389 2144 5397 2208
rect 5077 2128 5397 2144
rect 11363 27776 11683 27792
rect 11363 27712 11371 27776
rect 11435 27712 11451 27776
rect 11515 27712 11531 27776
rect 11595 27712 11611 27776
rect 11675 27712 11683 27776
rect 11363 26688 11683 27712
rect 11363 26624 11371 26688
rect 11435 26624 11451 26688
rect 11515 26624 11531 26688
rect 11595 26624 11611 26688
rect 11675 26624 11683 26688
rect 11363 25600 11683 26624
rect 11363 25536 11371 25600
rect 11435 25536 11451 25600
rect 11515 25536 11531 25600
rect 11595 25536 11611 25600
rect 11675 25536 11683 25600
rect 11363 24666 11683 25536
rect 11363 24512 11405 24666
rect 11641 24512 11683 24666
rect 11363 24448 11371 24512
rect 11675 24448 11683 24512
rect 11363 24430 11405 24448
rect 11641 24430 11683 24448
rect 11363 23424 11683 24430
rect 11363 23360 11371 23424
rect 11435 23360 11451 23424
rect 11515 23360 11531 23424
rect 11595 23360 11611 23424
rect 11675 23360 11683 23424
rect 11363 22336 11683 23360
rect 11363 22272 11371 22336
rect 11435 22272 11451 22336
rect 11515 22272 11531 22336
rect 11595 22272 11611 22336
rect 11675 22272 11683 22336
rect 11363 21248 11683 22272
rect 11363 21184 11371 21248
rect 11435 21184 11451 21248
rect 11515 21184 11531 21248
rect 11595 21184 11611 21248
rect 11675 21184 11683 21248
rect 11363 20160 11683 21184
rect 11363 20096 11371 20160
rect 11435 20096 11451 20160
rect 11515 20096 11531 20160
rect 11595 20096 11611 20160
rect 11675 20096 11683 20160
rect 11363 19072 11683 20096
rect 11363 19008 11371 19072
rect 11435 19008 11451 19072
rect 11515 19008 11531 19072
rect 11595 19008 11611 19072
rect 11675 19008 11683 19072
rect 11363 18274 11683 19008
rect 11363 18038 11405 18274
rect 11641 18038 11683 18274
rect 11363 17984 11683 18038
rect 11363 17920 11371 17984
rect 11435 17920 11451 17984
rect 11515 17920 11531 17984
rect 11595 17920 11611 17984
rect 11675 17920 11683 17984
rect 11363 16896 11683 17920
rect 11363 16832 11371 16896
rect 11435 16832 11451 16896
rect 11515 16832 11531 16896
rect 11595 16832 11611 16896
rect 11675 16832 11683 16896
rect 11363 15808 11683 16832
rect 11363 15744 11371 15808
rect 11435 15744 11451 15808
rect 11515 15744 11531 15808
rect 11595 15744 11611 15808
rect 11675 15744 11683 15808
rect 11363 14720 11683 15744
rect 11363 14656 11371 14720
rect 11435 14656 11451 14720
rect 11515 14656 11531 14720
rect 11595 14656 11611 14720
rect 11675 14656 11683 14720
rect 11363 13632 11683 14656
rect 11363 13568 11371 13632
rect 11435 13568 11451 13632
rect 11515 13568 11531 13632
rect 11595 13568 11611 13632
rect 11675 13568 11683 13632
rect 11363 12544 11683 13568
rect 11363 12480 11371 12544
rect 11435 12480 11451 12544
rect 11515 12480 11531 12544
rect 11595 12480 11611 12544
rect 11675 12480 11683 12544
rect 11363 11882 11683 12480
rect 11363 11646 11405 11882
rect 11641 11646 11683 11882
rect 11363 11456 11683 11646
rect 11363 11392 11371 11456
rect 11435 11392 11451 11456
rect 11515 11392 11531 11456
rect 11595 11392 11611 11456
rect 11675 11392 11683 11456
rect 11363 10368 11683 11392
rect 11363 10304 11371 10368
rect 11435 10304 11451 10368
rect 11515 10304 11531 10368
rect 11595 10304 11611 10368
rect 11675 10304 11683 10368
rect 11363 9280 11683 10304
rect 11363 9216 11371 9280
rect 11435 9216 11451 9280
rect 11515 9216 11531 9280
rect 11595 9216 11611 9280
rect 11675 9216 11683 9280
rect 11363 8192 11683 9216
rect 11363 8128 11371 8192
rect 11435 8128 11451 8192
rect 11515 8128 11531 8192
rect 11595 8128 11611 8192
rect 11675 8128 11683 8192
rect 11363 7104 11683 8128
rect 11363 7040 11371 7104
rect 11435 7040 11451 7104
rect 11515 7040 11531 7104
rect 11595 7040 11611 7104
rect 11675 7040 11683 7104
rect 11363 6016 11683 7040
rect 11363 5952 11371 6016
rect 11435 5952 11451 6016
rect 11515 5952 11531 6016
rect 11595 5952 11611 6016
rect 11675 5952 11683 6016
rect 11363 5490 11683 5952
rect 11363 5254 11405 5490
rect 11641 5254 11683 5490
rect 11363 4928 11683 5254
rect 11363 4864 11371 4928
rect 11435 4864 11451 4928
rect 11515 4864 11531 4928
rect 11595 4864 11611 4928
rect 11675 4864 11683 4928
rect 11363 3840 11683 4864
rect 11363 3776 11371 3840
rect 11435 3776 11451 3840
rect 11515 3776 11531 3840
rect 11595 3776 11611 3840
rect 11675 3776 11683 3840
rect 11363 2752 11683 3776
rect 11363 2688 11371 2752
rect 11435 2688 11451 2752
rect 11515 2688 11531 2752
rect 11595 2688 11611 2752
rect 11675 2688 11683 2752
rect 11363 2128 11683 2688
rect 12023 27232 12343 27792
rect 12023 27168 12031 27232
rect 12095 27168 12111 27232
rect 12175 27168 12191 27232
rect 12255 27168 12271 27232
rect 12335 27168 12343 27232
rect 12023 26144 12343 27168
rect 12023 26080 12031 26144
rect 12095 26080 12111 26144
rect 12175 26080 12191 26144
rect 12255 26080 12271 26144
rect 12335 26080 12343 26144
rect 12023 25326 12343 26080
rect 12023 25090 12065 25326
rect 12301 25090 12343 25326
rect 12023 25056 12343 25090
rect 12023 24992 12031 25056
rect 12095 24992 12111 25056
rect 12175 24992 12191 25056
rect 12255 24992 12271 25056
rect 12335 24992 12343 25056
rect 12023 23968 12343 24992
rect 12023 23904 12031 23968
rect 12095 23904 12111 23968
rect 12175 23904 12191 23968
rect 12255 23904 12271 23968
rect 12335 23904 12343 23968
rect 12023 22880 12343 23904
rect 12023 22816 12031 22880
rect 12095 22816 12111 22880
rect 12175 22816 12191 22880
rect 12255 22816 12271 22880
rect 12335 22816 12343 22880
rect 12023 21792 12343 22816
rect 12023 21728 12031 21792
rect 12095 21728 12111 21792
rect 12175 21728 12191 21792
rect 12255 21728 12271 21792
rect 12335 21728 12343 21792
rect 12023 20704 12343 21728
rect 12023 20640 12031 20704
rect 12095 20640 12111 20704
rect 12175 20640 12191 20704
rect 12255 20640 12271 20704
rect 12335 20640 12343 20704
rect 12023 19616 12343 20640
rect 12023 19552 12031 19616
rect 12095 19552 12111 19616
rect 12175 19552 12191 19616
rect 12255 19552 12271 19616
rect 12335 19552 12343 19616
rect 12023 18934 12343 19552
rect 12023 18698 12065 18934
rect 12301 18698 12343 18934
rect 12023 18528 12343 18698
rect 12023 18464 12031 18528
rect 12095 18464 12111 18528
rect 12175 18464 12191 18528
rect 12255 18464 12271 18528
rect 12335 18464 12343 18528
rect 12023 17440 12343 18464
rect 12023 17376 12031 17440
rect 12095 17376 12111 17440
rect 12175 17376 12191 17440
rect 12255 17376 12271 17440
rect 12335 17376 12343 17440
rect 12023 16352 12343 17376
rect 12023 16288 12031 16352
rect 12095 16288 12111 16352
rect 12175 16288 12191 16352
rect 12255 16288 12271 16352
rect 12335 16288 12343 16352
rect 12023 15264 12343 16288
rect 12023 15200 12031 15264
rect 12095 15200 12111 15264
rect 12175 15200 12191 15264
rect 12255 15200 12271 15264
rect 12335 15200 12343 15264
rect 12023 14176 12343 15200
rect 12023 14112 12031 14176
rect 12095 14112 12111 14176
rect 12175 14112 12191 14176
rect 12255 14112 12271 14176
rect 12335 14112 12343 14176
rect 12023 13088 12343 14112
rect 12023 13024 12031 13088
rect 12095 13024 12111 13088
rect 12175 13024 12191 13088
rect 12255 13024 12271 13088
rect 12335 13024 12343 13088
rect 12023 12542 12343 13024
rect 12023 12306 12065 12542
rect 12301 12306 12343 12542
rect 12023 12000 12343 12306
rect 12023 11936 12031 12000
rect 12095 11936 12111 12000
rect 12175 11936 12191 12000
rect 12255 11936 12271 12000
rect 12335 11936 12343 12000
rect 12023 10912 12343 11936
rect 12023 10848 12031 10912
rect 12095 10848 12111 10912
rect 12175 10848 12191 10912
rect 12255 10848 12271 10912
rect 12335 10848 12343 10912
rect 12023 9824 12343 10848
rect 12023 9760 12031 9824
rect 12095 9760 12111 9824
rect 12175 9760 12191 9824
rect 12255 9760 12271 9824
rect 12335 9760 12343 9824
rect 12023 8736 12343 9760
rect 12023 8672 12031 8736
rect 12095 8672 12111 8736
rect 12175 8672 12191 8736
rect 12255 8672 12271 8736
rect 12335 8672 12343 8736
rect 12023 7648 12343 8672
rect 12023 7584 12031 7648
rect 12095 7584 12111 7648
rect 12175 7584 12191 7648
rect 12255 7584 12271 7648
rect 12335 7584 12343 7648
rect 12023 6560 12343 7584
rect 12023 6496 12031 6560
rect 12095 6496 12111 6560
rect 12175 6496 12191 6560
rect 12255 6496 12271 6560
rect 12335 6496 12343 6560
rect 12023 6150 12343 6496
rect 12023 5914 12065 6150
rect 12301 5914 12343 6150
rect 12023 5472 12343 5914
rect 12023 5408 12031 5472
rect 12095 5408 12111 5472
rect 12175 5408 12191 5472
rect 12255 5408 12271 5472
rect 12335 5408 12343 5472
rect 12023 4384 12343 5408
rect 12023 4320 12031 4384
rect 12095 4320 12111 4384
rect 12175 4320 12191 4384
rect 12255 4320 12271 4384
rect 12335 4320 12343 4384
rect 12023 3296 12343 4320
rect 12023 3232 12031 3296
rect 12095 3232 12111 3296
rect 12175 3232 12191 3296
rect 12255 3232 12271 3296
rect 12335 3232 12343 3296
rect 12023 2208 12343 3232
rect 12023 2144 12031 2208
rect 12095 2144 12111 2208
rect 12175 2144 12191 2208
rect 12255 2144 12271 2208
rect 12335 2144 12343 2208
rect 12023 2128 12343 2144
rect 18309 27776 18629 27792
rect 18309 27712 18317 27776
rect 18381 27712 18397 27776
rect 18461 27712 18477 27776
rect 18541 27712 18557 27776
rect 18621 27712 18629 27776
rect 18309 26688 18629 27712
rect 18309 26624 18317 26688
rect 18381 26624 18397 26688
rect 18461 26624 18477 26688
rect 18541 26624 18557 26688
rect 18621 26624 18629 26688
rect 18309 25600 18629 26624
rect 18309 25536 18317 25600
rect 18381 25536 18397 25600
rect 18461 25536 18477 25600
rect 18541 25536 18557 25600
rect 18621 25536 18629 25600
rect 18309 24666 18629 25536
rect 18309 24512 18351 24666
rect 18587 24512 18629 24666
rect 18309 24448 18317 24512
rect 18621 24448 18629 24512
rect 18309 24430 18351 24448
rect 18587 24430 18629 24448
rect 18309 23424 18629 24430
rect 18309 23360 18317 23424
rect 18381 23360 18397 23424
rect 18461 23360 18477 23424
rect 18541 23360 18557 23424
rect 18621 23360 18629 23424
rect 18309 22336 18629 23360
rect 18309 22272 18317 22336
rect 18381 22272 18397 22336
rect 18461 22272 18477 22336
rect 18541 22272 18557 22336
rect 18621 22272 18629 22336
rect 18309 21248 18629 22272
rect 18309 21184 18317 21248
rect 18381 21184 18397 21248
rect 18461 21184 18477 21248
rect 18541 21184 18557 21248
rect 18621 21184 18629 21248
rect 18309 20160 18629 21184
rect 18309 20096 18317 20160
rect 18381 20096 18397 20160
rect 18461 20096 18477 20160
rect 18541 20096 18557 20160
rect 18621 20096 18629 20160
rect 18309 19072 18629 20096
rect 18309 19008 18317 19072
rect 18381 19008 18397 19072
rect 18461 19008 18477 19072
rect 18541 19008 18557 19072
rect 18621 19008 18629 19072
rect 18309 18274 18629 19008
rect 18309 18038 18351 18274
rect 18587 18038 18629 18274
rect 18309 17984 18629 18038
rect 18309 17920 18317 17984
rect 18381 17920 18397 17984
rect 18461 17920 18477 17984
rect 18541 17920 18557 17984
rect 18621 17920 18629 17984
rect 18309 16896 18629 17920
rect 18309 16832 18317 16896
rect 18381 16832 18397 16896
rect 18461 16832 18477 16896
rect 18541 16832 18557 16896
rect 18621 16832 18629 16896
rect 18309 15808 18629 16832
rect 18309 15744 18317 15808
rect 18381 15744 18397 15808
rect 18461 15744 18477 15808
rect 18541 15744 18557 15808
rect 18621 15744 18629 15808
rect 18309 14720 18629 15744
rect 18309 14656 18317 14720
rect 18381 14656 18397 14720
rect 18461 14656 18477 14720
rect 18541 14656 18557 14720
rect 18621 14656 18629 14720
rect 18309 13632 18629 14656
rect 18309 13568 18317 13632
rect 18381 13568 18397 13632
rect 18461 13568 18477 13632
rect 18541 13568 18557 13632
rect 18621 13568 18629 13632
rect 18309 12544 18629 13568
rect 18309 12480 18317 12544
rect 18381 12480 18397 12544
rect 18461 12480 18477 12544
rect 18541 12480 18557 12544
rect 18621 12480 18629 12544
rect 18309 11882 18629 12480
rect 18309 11646 18351 11882
rect 18587 11646 18629 11882
rect 18309 11456 18629 11646
rect 18309 11392 18317 11456
rect 18381 11392 18397 11456
rect 18461 11392 18477 11456
rect 18541 11392 18557 11456
rect 18621 11392 18629 11456
rect 18309 10368 18629 11392
rect 18309 10304 18317 10368
rect 18381 10304 18397 10368
rect 18461 10304 18477 10368
rect 18541 10304 18557 10368
rect 18621 10304 18629 10368
rect 18309 9280 18629 10304
rect 18309 9216 18317 9280
rect 18381 9216 18397 9280
rect 18461 9216 18477 9280
rect 18541 9216 18557 9280
rect 18621 9216 18629 9280
rect 18309 8192 18629 9216
rect 18309 8128 18317 8192
rect 18381 8128 18397 8192
rect 18461 8128 18477 8192
rect 18541 8128 18557 8192
rect 18621 8128 18629 8192
rect 18309 7104 18629 8128
rect 18309 7040 18317 7104
rect 18381 7040 18397 7104
rect 18461 7040 18477 7104
rect 18541 7040 18557 7104
rect 18621 7040 18629 7104
rect 18309 6016 18629 7040
rect 18309 5952 18317 6016
rect 18381 5952 18397 6016
rect 18461 5952 18477 6016
rect 18541 5952 18557 6016
rect 18621 5952 18629 6016
rect 18309 5490 18629 5952
rect 18309 5254 18351 5490
rect 18587 5254 18629 5490
rect 18309 4928 18629 5254
rect 18309 4864 18317 4928
rect 18381 4864 18397 4928
rect 18461 4864 18477 4928
rect 18541 4864 18557 4928
rect 18621 4864 18629 4928
rect 18309 3840 18629 4864
rect 18309 3776 18317 3840
rect 18381 3776 18397 3840
rect 18461 3776 18477 3840
rect 18541 3776 18557 3840
rect 18621 3776 18629 3840
rect 18309 2752 18629 3776
rect 18309 2688 18317 2752
rect 18381 2688 18397 2752
rect 18461 2688 18477 2752
rect 18541 2688 18557 2752
rect 18621 2688 18629 2752
rect 18309 2128 18629 2688
rect 18969 27232 19289 27792
rect 18969 27168 18977 27232
rect 19041 27168 19057 27232
rect 19121 27168 19137 27232
rect 19201 27168 19217 27232
rect 19281 27168 19289 27232
rect 18969 26144 19289 27168
rect 18969 26080 18977 26144
rect 19041 26080 19057 26144
rect 19121 26080 19137 26144
rect 19201 26080 19217 26144
rect 19281 26080 19289 26144
rect 18969 25326 19289 26080
rect 18969 25090 19011 25326
rect 19247 25090 19289 25326
rect 18969 25056 19289 25090
rect 18969 24992 18977 25056
rect 19041 24992 19057 25056
rect 19121 24992 19137 25056
rect 19201 24992 19217 25056
rect 19281 24992 19289 25056
rect 18969 23968 19289 24992
rect 18969 23904 18977 23968
rect 19041 23904 19057 23968
rect 19121 23904 19137 23968
rect 19201 23904 19217 23968
rect 19281 23904 19289 23968
rect 18969 22880 19289 23904
rect 18969 22816 18977 22880
rect 19041 22816 19057 22880
rect 19121 22816 19137 22880
rect 19201 22816 19217 22880
rect 19281 22816 19289 22880
rect 18969 21792 19289 22816
rect 18969 21728 18977 21792
rect 19041 21728 19057 21792
rect 19121 21728 19137 21792
rect 19201 21728 19217 21792
rect 19281 21728 19289 21792
rect 18969 20704 19289 21728
rect 18969 20640 18977 20704
rect 19041 20640 19057 20704
rect 19121 20640 19137 20704
rect 19201 20640 19217 20704
rect 19281 20640 19289 20704
rect 18969 19616 19289 20640
rect 18969 19552 18977 19616
rect 19041 19552 19057 19616
rect 19121 19552 19137 19616
rect 19201 19552 19217 19616
rect 19281 19552 19289 19616
rect 18969 18934 19289 19552
rect 18969 18698 19011 18934
rect 19247 18698 19289 18934
rect 18969 18528 19289 18698
rect 18969 18464 18977 18528
rect 19041 18464 19057 18528
rect 19121 18464 19137 18528
rect 19201 18464 19217 18528
rect 19281 18464 19289 18528
rect 18969 17440 19289 18464
rect 18969 17376 18977 17440
rect 19041 17376 19057 17440
rect 19121 17376 19137 17440
rect 19201 17376 19217 17440
rect 19281 17376 19289 17440
rect 18969 16352 19289 17376
rect 18969 16288 18977 16352
rect 19041 16288 19057 16352
rect 19121 16288 19137 16352
rect 19201 16288 19217 16352
rect 19281 16288 19289 16352
rect 18969 15264 19289 16288
rect 25255 27776 25575 27792
rect 25255 27712 25263 27776
rect 25327 27712 25343 27776
rect 25407 27712 25423 27776
rect 25487 27712 25503 27776
rect 25567 27712 25575 27776
rect 25255 26688 25575 27712
rect 25255 26624 25263 26688
rect 25327 26624 25343 26688
rect 25407 26624 25423 26688
rect 25487 26624 25503 26688
rect 25567 26624 25575 26688
rect 25255 25600 25575 26624
rect 25255 25536 25263 25600
rect 25327 25536 25343 25600
rect 25407 25536 25423 25600
rect 25487 25536 25503 25600
rect 25567 25536 25575 25600
rect 25255 24666 25575 25536
rect 25255 24512 25297 24666
rect 25533 24512 25575 24666
rect 25255 24448 25263 24512
rect 25567 24448 25575 24512
rect 25255 24430 25297 24448
rect 25533 24430 25575 24448
rect 25255 23424 25575 24430
rect 25255 23360 25263 23424
rect 25327 23360 25343 23424
rect 25407 23360 25423 23424
rect 25487 23360 25503 23424
rect 25567 23360 25575 23424
rect 25255 22336 25575 23360
rect 25255 22272 25263 22336
rect 25327 22272 25343 22336
rect 25407 22272 25423 22336
rect 25487 22272 25503 22336
rect 25567 22272 25575 22336
rect 25255 21248 25575 22272
rect 25255 21184 25263 21248
rect 25327 21184 25343 21248
rect 25407 21184 25423 21248
rect 25487 21184 25503 21248
rect 25567 21184 25575 21248
rect 25255 20160 25575 21184
rect 25255 20096 25263 20160
rect 25327 20096 25343 20160
rect 25407 20096 25423 20160
rect 25487 20096 25503 20160
rect 25567 20096 25575 20160
rect 25255 19072 25575 20096
rect 25255 19008 25263 19072
rect 25327 19008 25343 19072
rect 25407 19008 25423 19072
rect 25487 19008 25503 19072
rect 25567 19008 25575 19072
rect 25255 18274 25575 19008
rect 25255 18038 25297 18274
rect 25533 18038 25575 18274
rect 25255 17984 25575 18038
rect 25255 17920 25263 17984
rect 25327 17920 25343 17984
rect 25407 17920 25423 17984
rect 25487 17920 25503 17984
rect 25567 17920 25575 17984
rect 25255 16896 25575 17920
rect 25255 16832 25263 16896
rect 25327 16832 25343 16896
rect 25407 16832 25423 16896
rect 25487 16832 25503 16896
rect 25567 16832 25575 16896
rect 25255 15808 25575 16832
rect 25255 15744 25263 15808
rect 25327 15744 25343 15808
rect 25407 15744 25423 15808
rect 25487 15744 25503 15808
rect 25567 15744 25575 15808
rect 24899 15740 24965 15741
rect 24899 15676 24900 15740
rect 24964 15676 24965 15740
rect 24899 15675 24965 15676
rect 18969 15200 18977 15264
rect 19041 15200 19057 15264
rect 19121 15200 19137 15264
rect 19201 15200 19217 15264
rect 19281 15200 19289 15264
rect 18969 14176 19289 15200
rect 18969 14112 18977 14176
rect 19041 14112 19057 14176
rect 19121 14112 19137 14176
rect 19201 14112 19217 14176
rect 19281 14112 19289 14176
rect 18969 13088 19289 14112
rect 18969 13024 18977 13088
rect 19041 13024 19057 13088
rect 19121 13024 19137 13088
rect 19201 13024 19217 13088
rect 19281 13024 19289 13088
rect 18969 12542 19289 13024
rect 18969 12306 19011 12542
rect 19247 12306 19289 12542
rect 18969 12000 19289 12306
rect 18969 11936 18977 12000
rect 19041 11936 19057 12000
rect 19121 11936 19137 12000
rect 19201 11936 19217 12000
rect 19281 11936 19289 12000
rect 18969 10912 19289 11936
rect 18969 10848 18977 10912
rect 19041 10848 19057 10912
rect 19121 10848 19137 10912
rect 19201 10848 19217 10912
rect 19281 10848 19289 10912
rect 18969 9824 19289 10848
rect 18969 9760 18977 9824
rect 19041 9760 19057 9824
rect 19121 9760 19137 9824
rect 19201 9760 19217 9824
rect 19281 9760 19289 9824
rect 18969 8736 19289 9760
rect 18969 8672 18977 8736
rect 19041 8672 19057 8736
rect 19121 8672 19137 8736
rect 19201 8672 19217 8736
rect 19281 8672 19289 8736
rect 18969 7648 19289 8672
rect 24902 8261 24962 15675
rect 25255 14720 25575 15744
rect 25255 14656 25263 14720
rect 25327 14656 25343 14720
rect 25407 14656 25423 14720
rect 25487 14656 25503 14720
rect 25567 14656 25575 14720
rect 25255 13632 25575 14656
rect 25255 13568 25263 13632
rect 25327 13568 25343 13632
rect 25407 13568 25423 13632
rect 25487 13568 25503 13632
rect 25567 13568 25575 13632
rect 25255 12544 25575 13568
rect 25255 12480 25263 12544
rect 25327 12480 25343 12544
rect 25407 12480 25423 12544
rect 25487 12480 25503 12544
rect 25567 12480 25575 12544
rect 25255 11882 25575 12480
rect 25255 11646 25297 11882
rect 25533 11646 25575 11882
rect 25255 11456 25575 11646
rect 25255 11392 25263 11456
rect 25327 11392 25343 11456
rect 25407 11392 25423 11456
rect 25487 11392 25503 11456
rect 25567 11392 25575 11456
rect 25255 10368 25575 11392
rect 25255 10304 25263 10368
rect 25327 10304 25343 10368
rect 25407 10304 25423 10368
rect 25487 10304 25503 10368
rect 25567 10304 25575 10368
rect 25255 9280 25575 10304
rect 25255 9216 25263 9280
rect 25327 9216 25343 9280
rect 25407 9216 25423 9280
rect 25487 9216 25503 9280
rect 25567 9216 25575 9280
rect 24899 8260 24965 8261
rect 24899 8196 24900 8260
rect 24964 8196 24965 8260
rect 24899 8195 24965 8196
rect 18969 7584 18977 7648
rect 19041 7584 19057 7648
rect 19121 7584 19137 7648
rect 19201 7584 19217 7648
rect 19281 7584 19289 7648
rect 18969 6560 19289 7584
rect 18969 6496 18977 6560
rect 19041 6496 19057 6560
rect 19121 6496 19137 6560
rect 19201 6496 19217 6560
rect 19281 6496 19289 6560
rect 18969 6150 19289 6496
rect 18969 5914 19011 6150
rect 19247 5914 19289 6150
rect 18969 5472 19289 5914
rect 18969 5408 18977 5472
rect 19041 5408 19057 5472
rect 19121 5408 19137 5472
rect 19201 5408 19217 5472
rect 19281 5408 19289 5472
rect 18969 4384 19289 5408
rect 18969 4320 18977 4384
rect 19041 4320 19057 4384
rect 19121 4320 19137 4384
rect 19201 4320 19217 4384
rect 19281 4320 19289 4384
rect 18969 3296 19289 4320
rect 18969 3232 18977 3296
rect 19041 3232 19057 3296
rect 19121 3232 19137 3296
rect 19201 3232 19217 3296
rect 19281 3232 19289 3296
rect 18969 2208 19289 3232
rect 18969 2144 18977 2208
rect 19041 2144 19057 2208
rect 19121 2144 19137 2208
rect 19201 2144 19217 2208
rect 19281 2144 19289 2208
rect 18969 2128 19289 2144
rect 25255 8192 25575 9216
rect 25255 8128 25263 8192
rect 25327 8128 25343 8192
rect 25407 8128 25423 8192
rect 25487 8128 25503 8192
rect 25567 8128 25575 8192
rect 25255 7104 25575 8128
rect 25255 7040 25263 7104
rect 25327 7040 25343 7104
rect 25407 7040 25423 7104
rect 25487 7040 25503 7104
rect 25567 7040 25575 7104
rect 25255 6016 25575 7040
rect 25255 5952 25263 6016
rect 25327 5952 25343 6016
rect 25407 5952 25423 6016
rect 25487 5952 25503 6016
rect 25567 5952 25575 6016
rect 25255 5490 25575 5952
rect 25255 5254 25297 5490
rect 25533 5254 25575 5490
rect 25255 4928 25575 5254
rect 25255 4864 25263 4928
rect 25327 4864 25343 4928
rect 25407 4864 25423 4928
rect 25487 4864 25503 4928
rect 25567 4864 25575 4928
rect 25255 3840 25575 4864
rect 25255 3776 25263 3840
rect 25327 3776 25343 3840
rect 25407 3776 25423 3840
rect 25487 3776 25503 3840
rect 25567 3776 25575 3840
rect 25255 2752 25575 3776
rect 25255 2688 25263 2752
rect 25327 2688 25343 2752
rect 25407 2688 25423 2752
rect 25487 2688 25503 2752
rect 25567 2688 25575 2752
rect 25255 2128 25575 2688
rect 25915 27232 26235 27792
rect 25915 27168 25923 27232
rect 25987 27168 26003 27232
rect 26067 27168 26083 27232
rect 26147 27168 26163 27232
rect 26227 27168 26235 27232
rect 25915 26144 26235 27168
rect 25915 26080 25923 26144
rect 25987 26080 26003 26144
rect 26067 26080 26083 26144
rect 26147 26080 26163 26144
rect 26227 26080 26235 26144
rect 25915 25326 26235 26080
rect 25915 25090 25957 25326
rect 26193 25090 26235 25326
rect 25915 25056 26235 25090
rect 25915 24992 25923 25056
rect 25987 24992 26003 25056
rect 26067 24992 26083 25056
rect 26147 24992 26163 25056
rect 26227 24992 26235 25056
rect 25915 23968 26235 24992
rect 25915 23904 25923 23968
rect 25987 23904 26003 23968
rect 26067 23904 26083 23968
rect 26147 23904 26163 23968
rect 26227 23904 26235 23968
rect 25915 22880 26235 23904
rect 25915 22816 25923 22880
rect 25987 22816 26003 22880
rect 26067 22816 26083 22880
rect 26147 22816 26163 22880
rect 26227 22816 26235 22880
rect 25915 21792 26235 22816
rect 25915 21728 25923 21792
rect 25987 21728 26003 21792
rect 26067 21728 26083 21792
rect 26147 21728 26163 21792
rect 26227 21728 26235 21792
rect 25915 20704 26235 21728
rect 25915 20640 25923 20704
rect 25987 20640 26003 20704
rect 26067 20640 26083 20704
rect 26147 20640 26163 20704
rect 26227 20640 26235 20704
rect 25915 19616 26235 20640
rect 25915 19552 25923 19616
rect 25987 19552 26003 19616
rect 26067 19552 26083 19616
rect 26147 19552 26163 19616
rect 26227 19552 26235 19616
rect 25915 18934 26235 19552
rect 25915 18698 25957 18934
rect 26193 18698 26235 18934
rect 25915 18528 26235 18698
rect 25915 18464 25923 18528
rect 25987 18464 26003 18528
rect 26067 18464 26083 18528
rect 26147 18464 26163 18528
rect 26227 18464 26235 18528
rect 25915 17440 26235 18464
rect 25915 17376 25923 17440
rect 25987 17376 26003 17440
rect 26067 17376 26083 17440
rect 26147 17376 26163 17440
rect 26227 17376 26235 17440
rect 25915 16352 26235 17376
rect 25915 16288 25923 16352
rect 25987 16288 26003 16352
rect 26067 16288 26083 16352
rect 26147 16288 26163 16352
rect 26227 16288 26235 16352
rect 25915 15264 26235 16288
rect 25915 15200 25923 15264
rect 25987 15200 26003 15264
rect 26067 15200 26083 15264
rect 26147 15200 26163 15264
rect 26227 15200 26235 15264
rect 25915 14176 26235 15200
rect 25915 14112 25923 14176
rect 25987 14112 26003 14176
rect 26067 14112 26083 14176
rect 26147 14112 26163 14176
rect 26227 14112 26235 14176
rect 25915 13088 26235 14112
rect 25915 13024 25923 13088
rect 25987 13024 26003 13088
rect 26067 13024 26083 13088
rect 26147 13024 26163 13088
rect 26227 13024 26235 13088
rect 25915 12542 26235 13024
rect 25915 12306 25957 12542
rect 26193 12306 26235 12542
rect 25915 12000 26235 12306
rect 25915 11936 25923 12000
rect 25987 11936 26003 12000
rect 26067 11936 26083 12000
rect 26147 11936 26163 12000
rect 26227 11936 26235 12000
rect 25915 10912 26235 11936
rect 25915 10848 25923 10912
rect 25987 10848 26003 10912
rect 26067 10848 26083 10912
rect 26147 10848 26163 10912
rect 26227 10848 26235 10912
rect 25915 9824 26235 10848
rect 25915 9760 25923 9824
rect 25987 9760 26003 9824
rect 26067 9760 26083 9824
rect 26147 9760 26163 9824
rect 26227 9760 26235 9824
rect 25915 8736 26235 9760
rect 25915 8672 25923 8736
rect 25987 8672 26003 8736
rect 26067 8672 26083 8736
rect 26147 8672 26163 8736
rect 26227 8672 26235 8736
rect 25915 7648 26235 8672
rect 25915 7584 25923 7648
rect 25987 7584 26003 7648
rect 26067 7584 26083 7648
rect 26147 7584 26163 7648
rect 26227 7584 26235 7648
rect 25915 6560 26235 7584
rect 25915 6496 25923 6560
rect 25987 6496 26003 6560
rect 26067 6496 26083 6560
rect 26147 6496 26163 6560
rect 26227 6496 26235 6560
rect 25915 6150 26235 6496
rect 25915 5914 25957 6150
rect 26193 5914 26235 6150
rect 25915 5472 26235 5914
rect 25915 5408 25923 5472
rect 25987 5408 26003 5472
rect 26067 5408 26083 5472
rect 26147 5408 26163 5472
rect 26227 5408 26235 5472
rect 25915 4384 26235 5408
rect 25915 4320 25923 4384
rect 25987 4320 26003 4384
rect 26067 4320 26083 4384
rect 26147 4320 26163 4384
rect 26227 4320 26235 4384
rect 25915 3296 26235 4320
rect 25915 3232 25923 3296
rect 25987 3232 26003 3296
rect 26067 3232 26083 3296
rect 26147 3232 26163 3296
rect 26227 3232 26235 3296
rect 25915 2208 26235 3232
rect 25915 2144 25923 2208
rect 25987 2144 26003 2208
rect 26067 2144 26083 2208
rect 26147 2144 26163 2208
rect 26227 2144 26235 2208
rect 25915 2128 26235 2144
<< via4 >>
rect 4459 24512 4695 24666
rect 4459 24448 4489 24512
rect 4489 24448 4505 24512
rect 4505 24448 4569 24512
rect 4569 24448 4585 24512
rect 4585 24448 4649 24512
rect 4649 24448 4665 24512
rect 4665 24448 4695 24512
rect 4459 24430 4695 24448
rect 4459 18038 4695 18274
rect 4459 11646 4695 11882
rect 4459 5254 4695 5490
rect 5119 25090 5355 25326
rect 5119 18698 5355 18934
rect 5119 12306 5355 12542
rect 5119 5914 5355 6150
rect 11405 24512 11641 24666
rect 11405 24448 11435 24512
rect 11435 24448 11451 24512
rect 11451 24448 11515 24512
rect 11515 24448 11531 24512
rect 11531 24448 11595 24512
rect 11595 24448 11611 24512
rect 11611 24448 11641 24512
rect 11405 24430 11641 24448
rect 11405 18038 11641 18274
rect 11405 11646 11641 11882
rect 11405 5254 11641 5490
rect 12065 25090 12301 25326
rect 12065 18698 12301 18934
rect 12065 12306 12301 12542
rect 12065 5914 12301 6150
rect 18351 24512 18587 24666
rect 18351 24448 18381 24512
rect 18381 24448 18397 24512
rect 18397 24448 18461 24512
rect 18461 24448 18477 24512
rect 18477 24448 18541 24512
rect 18541 24448 18557 24512
rect 18557 24448 18587 24512
rect 18351 24430 18587 24448
rect 18351 18038 18587 18274
rect 18351 11646 18587 11882
rect 18351 5254 18587 5490
rect 19011 25090 19247 25326
rect 19011 18698 19247 18934
rect 25297 24512 25533 24666
rect 25297 24448 25327 24512
rect 25327 24448 25343 24512
rect 25343 24448 25407 24512
rect 25407 24448 25423 24512
rect 25423 24448 25487 24512
rect 25487 24448 25503 24512
rect 25503 24448 25533 24512
rect 25297 24430 25533 24448
rect 25297 18038 25533 18274
rect 19011 12306 19247 12542
rect 25297 11646 25533 11882
rect 19011 5914 19247 6150
rect 25297 5254 25533 5490
rect 25957 25090 26193 25326
rect 25957 18698 26193 18934
rect 25957 12306 26193 12542
rect 25957 5914 26193 6150
<< metal5 >>
rect 1056 25326 28936 25368
rect 1056 25090 5119 25326
rect 5355 25090 12065 25326
rect 12301 25090 19011 25326
rect 19247 25090 25957 25326
rect 26193 25090 28936 25326
rect 1056 25048 28936 25090
rect 1056 24666 28936 24708
rect 1056 24430 4459 24666
rect 4695 24430 11405 24666
rect 11641 24430 18351 24666
rect 18587 24430 25297 24666
rect 25533 24430 28936 24666
rect 1056 24388 28936 24430
rect 1056 18934 28936 18976
rect 1056 18698 5119 18934
rect 5355 18698 12065 18934
rect 12301 18698 19011 18934
rect 19247 18698 25957 18934
rect 26193 18698 28936 18934
rect 1056 18656 28936 18698
rect 1056 18274 28936 18316
rect 1056 18038 4459 18274
rect 4695 18038 11405 18274
rect 11641 18038 18351 18274
rect 18587 18038 25297 18274
rect 25533 18038 28936 18274
rect 1056 17996 28936 18038
rect 1056 12542 28936 12584
rect 1056 12306 5119 12542
rect 5355 12306 12065 12542
rect 12301 12306 19011 12542
rect 19247 12306 25957 12542
rect 26193 12306 28936 12542
rect 1056 12264 28936 12306
rect 1056 11882 28936 11924
rect 1056 11646 4459 11882
rect 4695 11646 11405 11882
rect 11641 11646 18351 11882
rect 18587 11646 25297 11882
rect 25533 11646 28936 11882
rect 1056 11604 28936 11646
rect 1056 6150 28936 6192
rect 1056 5914 5119 6150
rect 5355 5914 12065 6150
rect 12301 5914 19011 6150
rect 19247 5914 25957 6150
rect 26193 5914 28936 6150
rect 1056 5872 28936 5914
rect 1056 5490 28936 5532
rect 1056 5254 4459 5490
rect 4695 5254 11405 5490
rect 11641 5254 18351 5490
rect 18587 5254 25297 5490
rect 25533 5254 28936 5490
rect 1056 5212 28936 5254
use sky130_fd_sc_hd__xnor2_1  _112_
timestamp 0
transform 1 0 17572 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _113_
timestamp 0
transform 1 0 18216 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _114_
timestamp 0
transform -1 0 19504 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _115_
timestamp 0
transform 1 0 15272 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _116_
timestamp 0
transform 1 0 13340 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _117_
timestamp 0
transform 1 0 16652 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _118_
timestamp 0
transform 1 0 18768 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 0
transform -1 0 24748 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_2  _120_
timestamp 0
transform -1 0 21712 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _121_
timestamp 0
transform 1 0 21804 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _122_
timestamp 0
transform 1 0 19228 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 0
transform 1 0 19412 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _124_
timestamp 0
transform 1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _125_
timestamp 0
transform -1 0 18676 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _126_
timestamp 0
transform 1 0 20056 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _127_
timestamp 0
transform 1 0 16468 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  _128_
timestamp 0
transform 1 0 19136 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _129_
timestamp 0
transform -1 0 22264 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _130_
timestamp 0
transform -1 0 22080 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _131_
timestamp 0
transform 1 0 19872 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _132_
timestamp 0
transform 1 0 20884 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _133_
timestamp 0
transform 1 0 20332 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _134_
timestamp 0
transform 1 0 21068 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 0
transform -1 0 21528 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _136_
timestamp 0
transform 1 0 23184 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _137_
timestamp 0
transform 1 0 23460 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _138_
timestamp 0
transform 1 0 19228 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _139_
timestamp 0
transform 1 0 19780 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _140_
timestamp 0
transform -1 0 24932 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _141_
timestamp 0
transform -1 0 21712 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _142_
timestamp 0
transform -1 0 22540 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _143_
timestamp 0
transform -1 0 21252 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _144_
timestamp 0
transform -1 0 20332 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _145_
timestamp 0
transform -1 0 24288 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _146_
timestamp 0
transform 1 0 21896 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _147_
timestamp 0
transform 1 0 22172 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _148_
timestamp 0
transform -1 0 22540 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _149_
timestamp 0
transform 1 0 24932 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _150_
timestamp 0
transform 1 0 22632 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _151_
timestamp 0
transform 1 0 22356 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _152_
timestamp 0
transform -1 0 23828 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _153_
timestamp 0
transform 1 0 23000 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _154_
timestamp 0
transform 1 0 22540 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _155_
timestamp 0
transform -1 0 21252 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _156_
timestamp 0
transform 1 0 21804 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _157_
timestamp 0
transform -1 0 20792 0 1 3264
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 0
transform 1 0 20240 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _159_
timestamp 0
transform 1 0 22724 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _160_
timestamp 0
transform -1 0 23276 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _161_
timestamp 0
transform -1 0 22724 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _162_
timestamp 0
transform -1 0 21988 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _163_
timestamp 0
transform -1 0 23092 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _164_
timestamp 0
transform 1 0 21804 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _165_
timestamp 0
transform -1 0 23736 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _166_
timestamp 0
transform -1 0 23184 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _167_
timestamp 0
transform 1 0 23736 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _168_
timestamp 0
transform -1 0 23644 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _169_
timestamp 0
transform -1 0 23368 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _170_
timestamp 0
transform 1 0 24748 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _171_
timestamp 0
transform 1 0 25116 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _172_
timestamp 0
transform 1 0 24104 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _173_
timestamp 0
transform -1 0 25760 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _174_
timestamp 0
transform -1 0 25116 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _175_
timestamp 0
transform 1 0 23368 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _176_
timestamp 0
transform -1 0 22816 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _177_
timestamp 0
transform 1 0 21988 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _178_
timestamp 0
transform 1 0 22816 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _179_
timestamp 0
transform -1 0 24104 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _180_
timestamp 0
transform 1 0 22264 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _181_
timestamp 0
transform 1 0 22632 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _182_
timestamp 0
transform -1 0 24012 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _183_
timestamp 0
transform 1 0 18676 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _184_
timestamp 0
transform 1 0 20332 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _185_
timestamp 0
transform 1 0 19320 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _186_
timestamp 0
transform 1 0 21068 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _187_
timestamp 0
transform -1 0 19412 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _188_
timestamp 0
transform 1 0 16284 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _189_
timestamp 0
transform 1 0 17664 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp 0
transform 1 0 18768 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _191_
timestamp 0
transform -1 0 17664 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _192_
timestamp 0
transform 1 0 17204 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _193_
timestamp 0
transform -1 0 18676 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _194_
timestamp 0
transform 1 0 17756 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _195_
timestamp 0
transform -1 0 20792 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 0
transform 1 0 19412 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _197_
timestamp 0
transform -1 0 20976 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _198_
timestamp 0
transform -1 0 21252 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _199_
timestamp 0
transform -1 0 21068 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _200_
timestamp 0
transform 1 0 18308 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _201_
timestamp 0
transform -1 0 18768 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _202_
timestamp 0
transform -1 0 18676 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _203_
timestamp 0
transform 1 0 17204 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _204_
timestamp 0
transform 1 0 17480 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _205_
timestamp 0
transform -1 0 20976 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _206_
timestamp 0
transform 1 0 19228 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _207_
timestamp 0
transform 1 0 20056 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _208_
timestamp 0
transform -1 0 18400 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _209_
timestamp 0
transform 1 0 18400 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _210_
timestamp 0
transform 1 0 17204 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _211_
timestamp 0
transform 1 0 17296 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _212_
timestamp 0
transform -1 0 14996 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _213_
timestamp 0
transform 1 0 14996 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _214_
timestamp 0
transform -1 0 14904 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _215_
timestamp 0
transform 1 0 14904 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _216_
timestamp 0
transform 1 0 16652 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _217_
timestamp 0
transform -1 0 16284 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _218_
timestamp 0
transform 1 0 14352 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _219_
timestamp 0
transform 1 0 14076 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _220_
timestamp 0
transform 1 0 15456 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _221_
timestamp 0
transform 1 0 14904 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _222_
timestamp 0
transform 1 0 16652 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _223_
timestamp 0
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _224_
timestamp 0
transform 1 0 18676 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _225_
timestamp 0
transform 1 0 19780 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _226_
timestamp 0
transform -1 0 22816 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _227_
timestamp 0
transform 1 0 22632 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _228_
timestamp 0
transform 1 0 23276 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _229_
timestamp 0
transform 1 0 22172 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _230_
timestamp 0
transform 1 0 19688 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _231_
timestamp 0
transform 1 0 21804 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _232_
timestamp 0
transform 1 0 19780 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _233_
timestamp 0
transform 1 0 24380 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _234_
timestamp 0
transform 1 0 24380 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _235_
timestamp 0
transform 1 0 24196 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _236_
timestamp 0
transform 1 0 20148 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _237_
timestamp 0
transform -1 0 21896 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _238_
timestamp 0
transform 1 0 23368 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _239_
timestamp 0
transform -1 0 20332 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _240_
timestamp 0
transform 1 0 17848 0 -1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _241_
timestamp 0
transform 1 0 15824 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _242_
timestamp 0
transform 1 0 16652 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _243_
timestamp 0
transform 1 0 16560 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _244_
timestamp 0
transform 1 0 16652 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _245_
timestamp 0
transform 1 0 19228 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _246_
timestamp 0
transform 1 0 18400 0 -1 7616
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _247_
timestamp 0
transform 1 0 16376 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _248_
timestamp 0
transform -1 0 20056 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _249_
timestamp 0
transform 1 0 16928 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _250_
timestamp 0
transform 1 0 16192 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _251_
timestamp 0
transform 1 0 14168 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _252_
timestamp 0
transform 1 0 14076 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _253_
timestamp 0
transform -1 0 16560 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _254_
timestamp 0
transform 1 0 13892 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _255_
timestamp 0
transform 1 0 14352 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _256_
timestamp 0
transform 1 0 15640 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 0
transform -1 0 21896 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 0
transform -1 0 17480 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 0
transform -1 0 17480 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 0
transform 1 0 20792 0 1 3264
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 0
transform 1 0 21896 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout13
timestamp 0
transform 1 0 18400 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout14
timestamp 0
transform -1 0 16468 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout15
timestamp 0
transform -1 0 21436 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  fanout16
timestamp 0
transform 1 0 18768 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_13
timestamp 0
transform 1 0 2300 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_25
timestamp 0
transform 1 0 3404 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 0
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 0
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_90
timestamp 0
transform 1 0 9384 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_102
timestamp 0
transform 1 0 10488 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_110
timestamp 0
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 0
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 0
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 0
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 0
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 0
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 0
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_181
timestamp 0
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_188
timestamp 0
transform 1 0 18400 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_197
timestamp 0
transform 1 0 19228 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_203
timestamp 0
transform 1 0 19780 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_207
timestamp 0
transform 1 0 20148 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_211
timestamp 0
transform 1 0 20516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 0
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_225
timestamp 0
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_241
timestamp 0
transform 1 0 23276 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 0
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 0
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 0
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 0
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_281
timestamp 0
transform 1 0 26956 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_286
timestamp 0
transform 1 0 27416 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_298
timestamp 0
transform 1 0 28520 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 0
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 0
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 0
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 0
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 0
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 0
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 0
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 0
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 0
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 0
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 0
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 0
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 0
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 0
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_169
timestamp 0
transform 1 0 16652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_178
timestamp 0
transform 1 0 17480 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 0
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_253
timestamp 0
transform 1 0 24380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_265
timestamp 0
transform 1 0 25484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_277
timestamp 0
transform 1 0 26588 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 0
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_293
timestamp 0
transform 1 0 28060 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 0
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 0
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 0
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 0
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 0
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 0
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 0
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 0
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 0
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 0
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 0
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_165
timestamp 0
transform 1 0 16284 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_194
timestamp 0
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 0
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 0
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_273
timestamp 0
transform 1 0 26220 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_285
timestamp 0
transform 1 0 27324 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_297
timestamp 0
transform 1 0 28428 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 0
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 0
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 0
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 0
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 0
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 0
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 0
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 0
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 0
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 0
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 0
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 0
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 0
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_161
timestamp 0
transform 1 0 15916 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_169
timestamp 0
transform 1 0 16652 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_185
timestamp 0
transform 1 0 18124 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_202
timestamp 0
transform 1 0 19688 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 0
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_254
timestamp 0
transform 1 0 24472 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_258
timestamp 0
transform 1 0 24840 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_267
timestamp 0
transform 1 0 25668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 0
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 0
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_293
timestamp 0
transform 1 0 28060 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 0
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 0
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 0
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 0
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 0
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 0
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 0
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 0
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 0
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 0
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 0
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_153
timestamp 0
transform 1 0 15180 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_159
timestamp 0
transform 1 0 15732 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_180
timestamp 0
transform 1 0 17664 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_220
timestamp 0
transform 1 0 21344 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_239
timestamp 0
transform 1 0 23092 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_246
timestamp 0
transform 1 0 23736 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_273
timestamp 0
transform 1 0 26220 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_285
timestamp 0
transform 1 0 27324 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_297
timestamp 0
transform 1 0 28428 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 0
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 0
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 0
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 0
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 0
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 0
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 0
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 0
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 0
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 0
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 0
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 0
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 0
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 0
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 0
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 0
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_222
timestamp 0
transform 1 0 21528 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_229
timestamp 0
transform 1 0 22172 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_236
timestamp 0
transform 1 0 22816 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_249
timestamp 0
transform 1 0 24012 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_260
timestamp 0
transform 1 0 25024 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_270
timestamp 0
transform 1 0 25944 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_278
timestamp 0
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 0
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_293
timestamp 0
transform 1 0 28060 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 0
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 0
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 0
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 0
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 0
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 0
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 0
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 0
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 0
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 0
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 0
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 0
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_153
timestamp 0
transform 1 0 15180 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_157
timestamp 0
transform 1 0 15548 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_205
timestamp 0
transform 1 0 19964 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_250
timestamp 0
transform 1 0 24104 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_267
timestamp 0
transform 1 0 25668 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_279
timestamp 0
transform 1 0 26772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_291
timestamp 0
transform 1 0 27876 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 0
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 0
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 0
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 0
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 0
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 0
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 0
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 0
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 0
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 0
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 0
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 0
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 0
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 0
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 0
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_212
timestamp 0
transform 1 0 20608 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_219
timestamp 0
transform 1 0 21252 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 0
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_225
timestamp 0
transform 1 0 21804 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_229
timestamp 0
transform 1 0 22172 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_235
timestamp 0
transform 1 0 22724 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_243
timestamp 0
transform 1 0 23460 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_250
timestamp 0
transform 1 0 24104 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_281
timestamp 0
transform 1 0 26956 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 0
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 0
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 0
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 0
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 0
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 0
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 0
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 0
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 0
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 0
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 0
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 0
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 0
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_165
timestamp 0
transform 1 0 16284 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_187
timestamp 0
transform 1 0 18308 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 0
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_197
timestamp 0
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_205
timestamp 0
transform 1 0 19964 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_249
timestamp 0
transform 1 0 24012 0 1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_268
timestamp 0
transform 1 0 25760 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_280
timestamp 0
transform 1 0 26864 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_292
timestamp 0
transform 1 0 27968 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_298
timestamp 0
transform 1 0 28520 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 0
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 0
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 0
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 0
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 0
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 0
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 0
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 0
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 0
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 0
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 0
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 0
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_137
timestamp 0
transform 1 0 13708 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_145
timestamp 0
transform 1 0 14444 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_169
timestamp 0
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_240
timestamp 0
transform 1 0 23184 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_262
timestamp 0
transform 1 0 25208 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_274
timestamp 0
transform 1 0 26312 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 0
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_293
timestamp 0
transform 1 0 28060 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 0
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 0
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 0
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 0
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 0
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 0
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 0
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 0
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 0
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 0
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 0
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 0
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 0
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_153
timestamp 0
transform 1 0 15180 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_157
timestamp 0
transform 1 0 15548 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_186
timestamp 0
transform 1 0 18216 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_263
timestamp 0
transform 1 0 25300 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_275
timestamp 0
transform 1 0 26404 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_287
timestamp 0
transform 1 0 27508 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 0
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 0
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 0
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 0
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 0
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 0
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 0
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 0
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 0
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 0
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 0
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_137
timestamp 0
transform 1 0 13708 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_159
timestamp 0
transform 1 0 15732 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 0
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_261
timestamp 0
transform 1 0 25116 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_273
timestamp 0
transform 1 0 26220 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 0
transform 1 0 26772 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 0
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_293
timestamp 0
transform 1 0 28060 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_6
timestamp 0
transform 1 0 1656 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_18
timestamp 0
transform 1 0 2760 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_26
timestamp 0
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 0
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 0
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 0
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 0
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 0
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 0
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 0
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 0
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 0
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 0
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_153
timestamp 0
transform 1 0 15180 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_165
timestamp 0
transform 1 0 16284 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_191
timestamp 0
transform 1 0 18676 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 0
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_197
timestamp 0
transform 1 0 19228 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_211
timestamp 0
transform 1 0 20516 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_247
timestamp 0
transform 1 0 23828 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 0
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_257
timestamp 0
transform 1 0 24748 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_269
timestamp 0
transform 1 0 25852 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_281
timestamp 0
transform 1 0 26956 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_293
timestamp 0
transform 1 0 28060 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 0
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 0
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 0
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 0
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 0
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 0
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 0
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 0
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 0
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 0
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 0
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 0
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_137
timestamp 0
transform 1 0 13708 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_153
timestamp 0
transform 1 0 15180 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 0
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 0
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_169
timestamp 0
transform 1 0 16652 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_191
timestamp 0
transform 1 0 18676 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_195
timestamp 0
transform 1 0 19044 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_219
timestamp 0
transform 1 0 21252 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 0
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_225
timestamp 0
transform 1 0 21804 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_246
timestamp 0
transform 1 0 23736 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_258
timestamp 0
transform 1 0 24840 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_270
timestamp 0
transform 1 0 25944 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_278
timestamp 0
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_281
timestamp 0
transform 1 0 26956 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_293
timestamp 0
transform 1 0 28060 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 0
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 0
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 0
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 0
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 0
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 0
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 0
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 0
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 0
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 0
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 0
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 0
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_169
timestamp 0
transform 1 0 16652 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_192
timestamp 0
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_197
timestamp 0
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_203
timestamp 0
transform 1 0 19780 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_212
timestamp 0
transform 1 0 20608 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_228
timestamp 0
transform 1 0 22080 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 0
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 0
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_277
timestamp 0
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_289
timestamp 0
transform 1 0 27692 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_297
timestamp 0
transform 1 0 28428 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 0
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 0
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 0
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 0
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 0
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 0
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 0
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 0
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 0
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 0
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 0
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 0
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_137
timestamp 0
transform 1 0 13708 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_141
timestamp 0
transform 1 0 14076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_162
timestamp 0
transform 1 0 16008 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_211
timestamp 0
transform 1 0 20516 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_222
timestamp 0
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_233
timestamp 0
transform 1 0 22540 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_257
timestamp 0
transform 1 0 24748 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_269
timestamp 0
transform 1 0 25852 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_277
timestamp 0
transform 1 0 26588 0 -1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_281
timestamp 0
transform 1 0 26956 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_293
timestamp 0
transform 1 0 28060 0 -1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 0
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 0
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 0
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 0
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 0
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 0
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 0
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 0
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 0
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 0
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_141
timestamp 0
transform 1 0 14076 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_162
timestamp 0
transform 1 0 16008 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_184
timestamp 0
transform 1 0 18032 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_214
timestamp 0
transform 1 0 20792 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_236
timestamp 0
transform 1 0 22816 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_248
timestamp 0
transform 1 0 23920 0 1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_253
timestamp 0
transform 1 0 24380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_265
timestamp 0
transform 1 0 25484 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_277
timestamp 0
transform 1 0 26588 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_289
timestamp 0
transform 1 0 27692 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_297
timestamp 0
transform 1 0 28428 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 0
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 0
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 0
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 0
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 0
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 0
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 0
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 0
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 0
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 0
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 0
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 0
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_137
timestamp 0
transform 1 0 13708 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_143
timestamp 0
transform 1 0 14260 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_164
timestamp 0
transform 1 0 16192 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_169
timestamp 0
transform 1 0 16652 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_202
timestamp 0
transform 1 0 19688 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 0
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_237
timestamp 0
transform 1 0 22908 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_249
timestamp 0
transform 1 0 24012 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_261
timestamp 0
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_273
timestamp 0
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 0
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_281
timestamp 0
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_293
timestamp 0
transform 1 0 28060 0 -1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 0
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 0
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 0
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 0
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 0
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 0
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 0
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 0
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 0
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 0
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 0
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 0
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_141
timestamp 0
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_149
timestamp 0
transform 1 0 14812 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_153
timestamp 0
transform 1 0 15180 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_157
timestamp 0
transform 1 0 15548 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_178
timestamp 0
transform 1 0 17480 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_186
timestamp 0
transform 1 0 18216 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_194
timestamp 0
transform 1 0 18952 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_197
timestamp 0
transform 1 0 19228 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_209
timestamp 0
transform 1 0 20332 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_221
timestamp 0
transform 1 0 21436 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_233
timestamp 0
transform 1 0 22540 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_245
timestamp 0
transform 1 0 23644 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 0
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_253
timestamp 0
transform 1 0 24380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_265
timestamp 0
transform 1 0 25484 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_277
timestamp 0
transform 1 0 26588 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_289
timestamp 0
transform 1 0 27692 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_297
timestamp 0
transform 1 0 28428 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_3
timestamp 0
transform 1 0 1380 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_15
timestamp 0
transform 1 0 2484 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_27
timestamp 0
transform 1 0 3588 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_39
timestamp 0
transform 1 0 4692 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_51
timestamp 0
transform 1 0 5796 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_55
timestamp 0
transform 1 0 6164 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 0
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 0
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 0
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 0
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 0
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 0
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 0
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 0
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_149
timestamp 0
transform 1 0 14812 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_155
timestamp 0
transform 1 0 15364 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_200
timestamp 0
transform 1 0 19504 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_212
timestamp 0
transform 1 0 20608 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_225
timestamp 0
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_237
timestamp 0
transform 1 0 22908 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_249
timestamp 0
transform 1 0 24012 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_261
timestamp 0
transform 1 0 25116 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_273
timestamp 0
transform 1 0 26220 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_279
timestamp 0
transform 1 0 26772 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 0
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_293
timestamp 0
transform 1 0 28060 0 -1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 0
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 0
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 0
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 0
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 0
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 0
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 0
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 0
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 0
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 0
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 0
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 0
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 0
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 0
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_153
timestamp 0
transform 1 0 15180 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_161
timestamp 0
transform 1 0 15916 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_170
timestamp 0
transform 1 0 16744 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_182
timestamp 0
transform 1 0 17848 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_194
timestamp 0
transform 1 0 18952 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_197
timestamp 0
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_209
timestamp 0
transform 1 0 20332 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_221
timestamp 0
transform 1 0 21436 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_233
timestamp 0
transform 1 0 22540 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_245
timestamp 0
transform 1 0 23644 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_251
timestamp 0
transform 1 0 24196 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_253
timestamp 0
transform 1 0 24380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_265
timestamp 0
transform 1 0 25484 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_277
timestamp 0
transform 1 0 26588 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_289
timestamp 0
transform 1 0 27692 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_297
timestamp 0
transform 1 0 28428 0 1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 0
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 0
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 0
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 0
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 0
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 0
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 0
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 0
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 0
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 0
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 0
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 0
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 0
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 0
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 0
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_149
timestamp 0
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 0
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 0
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 0
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_181
timestamp 0
transform 1 0 17756 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_193
timestamp 0
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_205
timestamp 0
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_217
timestamp 0
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 0
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_225
timestamp 0
transform 1 0 21804 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_237
timestamp 0
transform 1 0 22908 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_249
timestamp 0
transform 1 0 24012 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_261
timestamp 0
transform 1 0 25116 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_273
timestamp 0
transform 1 0 26220 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_279
timestamp 0
transform 1 0 26772 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_281
timestamp 0
transform 1 0 26956 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_293
timestamp 0
transform 1 0 28060 0 -1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 0
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 0
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 0
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 0
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 0
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 0
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 0
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 0
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 0
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 0
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 0
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 0
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 0
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 0
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 0
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 0
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 0
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 0
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_177
timestamp 0
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_189
timestamp 0
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 0
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 0
transform 1 0 19228 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_209
timestamp 0
transform 1 0 20332 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_221
timestamp 0
transform 1 0 21436 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_233
timestamp 0
transform 1 0 22540 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_245
timestamp 0
transform 1 0 23644 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 0
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 0
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 0
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 0
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_289
timestamp 0
transform 1 0 27692 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_297
timestamp 0
transform 1 0 28428 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 0
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 0
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 0
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 0
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 0
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 0
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 0
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 0
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 0
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 0
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 0
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 0
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 0
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 0
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 0
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 0
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 0
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 0
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 0
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_181
timestamp 0
transform 1 0 17756 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_193
timestamp 0
transform 1 0 18860 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_205
timestamp 0
transform 1 0 19964 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_217
timestamp 0
transform 1 0 21068 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 0
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_225
timestamp 0
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_237
timestamp 0
transform 1 0 22908 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_249
timestamp 0
transform 1 0 24012 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_261
timestamp 0
transform 1 0 25116 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_273
timestamp 0
transform 1 0 26220 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 0
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 0
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_293
timestamp 0
transform 1 0 28060 0 -1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 0
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 0
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 0
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 0
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 0
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 0
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 0
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 0
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 0
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 0
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 0
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 0
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 0
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 0
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 0
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 0
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 0
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_165
timestamp 0
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_177
timestamp 0
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_189
timestamp 0
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 0
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 0
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_209
timestamp 0
transform 1 0 20332 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_221
timestamp 0
transform 1 0 21436 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_233
timestamp 0
transform 1 0 22540 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_245
timestamp 0
transform 1 0 23644 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 0
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_253
timestamp 0
transform 1 0 24380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_265
timestamp 0
transform 1 0 25484 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_277
timestamp 0
transform 1 0 26588 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_289
timestamp 0
transform 1 0 27692 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_297
timestamp 0
transform 1 0 28428 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 0
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 0
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 0
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 0
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 0
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 0
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 0
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 0
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 0
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 0
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 0
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 0
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 0
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 0
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 0
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 0
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 0
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 0
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 0
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 0
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_193
timestamp 0
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 0
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 0
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 0
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_225
timestamp 0
transform 1 0 21804 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_237
timestamp 0
transform 1 0 22908 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_249
timestamp 0
transform 1 0 24012 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_261
timestamp 0
transform 1 0 25116 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_273
timestamp 0
transform 1 0 26220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_279
timestamp 0
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 0
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_293
timestamp 0
transform 1 0 28060 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 0
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 0
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 0
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 0
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 0
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 0
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 0
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 0
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 0
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 0
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 0
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 0
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 0
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 0
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 0
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 0
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 0
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 0
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 0
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_189
timestamp 0
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 0
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 0
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 0
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_221
timestamp 0
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_233
timestamp 0
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_245
timestamp 0
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 0
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 0
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_265
timestamp 0
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_277
timestamp 0
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_289
timestamp 0
transform 1 0 27692 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_297
timestamp 0
transform 1 0 28428 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 0
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 0
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 0
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 0
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 0
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 0
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 0
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 0
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 0
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 0
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 0
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 0
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 0
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 0
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 0
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 0
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 0
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 0
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 0
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_181
timestamp 0
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_193
timestamp 0
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_205
timestamp 0
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_217
timestamp 0
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 0
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 0
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_237
timestamp 0
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_249
timestamp 0
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_261
timestamp 0
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_273
timestamp 0
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 0
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 0
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_293
timestamp 0
transform 1 0 28060 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 0
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 0
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 0
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 0
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 0
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 0
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 0
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 0
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 0
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 0
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 0
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 0
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 0
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 0
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 0
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 0
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 0
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 0
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_177
timestamp 0
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 0
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 0
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 0
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 0
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_221
timestamp 0
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_233
timestamp 0
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_245
timestamp 0
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 0
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 0
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_265
timestamp 0
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_277
timestamp 0
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_289
timestamp 0
transform 1 0 27692 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_297
timestamp 0
transform 1 0 28428 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 0
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 0
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 0
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 0
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 0
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 0
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 0
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 0
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 0
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_93
timestamp 0
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 0
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 0
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 0
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 0
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 0
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 0
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 0
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 0
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 0
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 0
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_193
timestamp 0
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_205
timestamp 0
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_217
timestamp 0
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 0
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 0
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 0
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 0
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_261
timestamp 0
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_273
timestamp 0
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 0
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 0
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_293
timestamp 0
transform 1 0 28060 0 -1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_13
timestamp 0
transform 1 0 2300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_25
timestamp 0
transform 1 0 3404 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 0
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 0
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 0
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 0
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 0
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 0
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 0
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 0
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 0
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 0
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 0
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 0
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 0
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 0
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp 0
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_177
timestamp 0
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp 0
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 0
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 0
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_209
timestamp 0
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_221
timestamp 0
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_233
timestamp 0
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_245
timestamp 0
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 0
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 0
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 0
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 0
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_289
timestamp 0
transform 1 0 27692 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_297
timestamp 0
transform 1 0 28428 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 0
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 0
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 0
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 0
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 0
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 0
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 0
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 0
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 0
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 0
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 0
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 0
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 0
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 0
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 0
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 0
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 0
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 0
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 0
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_181
timestamp 0
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_193
timestamp 0
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_205
timestamp 0
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 0
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 0
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 0
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 0
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 0
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_261
timestamp 0
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_273
timestamp 0
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 0
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 0
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_293
timestamp 0
transform 1 0 28060 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 0
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 0
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 0
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 0
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 0
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 0
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 0
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 0
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 0
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 0
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 0
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 0
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 0
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 0
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 0
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 0
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 0
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_165
timestamp 0
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_177
timestamp 0
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_189
timestamp 0
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 0
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 0
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 0
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 0
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_233
timestamp 0
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 0
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 0
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 0
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 0
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_277
timestamp 0
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_289
timestamp 0
transform 1 0 27692 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_297
timestamp 0
transform 1 0 28428 0 1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 0
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 0
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 0
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 0
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 0
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 0
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 0
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 0
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 0
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_93
timestamp 0
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_105
timestamp 0
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 0
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 0
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 0
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_137
timestamp 0
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_149
timestamp 0
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_161
timestamp 0
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 0
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 0
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_181
timestamp 0
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_193
timestamp 0
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_205
timestamp 0
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_217
timestamp 0
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 0
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 0
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_237
timestamp 0
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_249
timestamp 0
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_261
timestamp 0
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_273
timestamp 0
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_279
timestamp 0
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 0
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_293
timestamp 0
transform 1 0 28060 0 -1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 0
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 0
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 0
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 0
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 0
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_53
timestamp 0
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_65
timestamp 0
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_77
timestamp 0
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 0
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 0
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_97
timestamp 0
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_109
timestamp 0
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_121
timestamp 0
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_133
timestamp 0
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 0
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 0
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_153
timestamp 0
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_165
timestamp 0
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_177
timestamp 0
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_189
timestamp 0
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 0
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_197
timestamp 0
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_209
timestamp 0
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_221
timestamp 0
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_233
timestamp 0
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_245
timestamp 0
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 0
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_253
timestamp 0
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_265
timestamp 0
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_277
timestamp 0
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_289
timestamp 0
transform 1 0 27692 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_297
timestamp 0
transform 1 0 28428 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 0
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 0
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 0
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_39
timestamp 0
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 0
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 0
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 0
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 0
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_81
timestamp 0
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_93
timestamp 0
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_105
timestamp 0
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 0
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 0
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_125
timestamp 0
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_137
timestamp 0
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_149
timestamp 0
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_161
timestamp 0
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 0
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 0
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_181
timestamp 0
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_193
timestamp 0
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_205
timestamp 0
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_217
timestamp 0
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 0
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 0
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_237
timestamp 0
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_249
timestamp 0
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_261
timestamp 0
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_273
timestamp 0
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_279
timestamp 0
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 0
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_293
timestamp 0
transform 1 0 28060 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 0
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 0
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 0
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 0
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 0
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_53
timestamp 0
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_65
timestamp 0
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_77
timestamp 0
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 0
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_85
timestamp 0
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_97
timestamp 0
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 0
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_121
timestamp 0
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 0
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 0
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_141
timestamp 0
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_153
timestamp 0
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_165
timestamp 0
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_177
timestamp 0
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_189
timestamp 0
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 0
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_197
timestamp 0
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_209
timestamp 0
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_221
timestamp 0
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_233
timestamp 0
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_245
timestamp 0
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 0
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 0
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_265
timestamp 0
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_277
timestamp 0
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_289
timestamp 0
transform 1 0 27692 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_297
timestamp 0
transform 1 0 28428 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 0
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 0
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 0
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 0
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 0
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 0
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 0
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 0
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_81
timestamp 0
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_93
timestamp 0
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_105
timestamp 0
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 0
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 0
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_125
timestamp 0
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_137
timestamp 0
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_149
timestamp 0
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_161
timestamp 0
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 0
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_169
timestamp 0
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_181
timestamp 0
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_193
timestamp 0
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_205
timestamp 0
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_217
timestamp 0
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 0
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_225
timestamp 0
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_237
timestamp 0
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_249
timestamp 0
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_261
timestamp 0
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_273
timestamp 0
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 0
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 0
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_293
timestamp 0
transform 1 0 28060 0 -1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 0
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 0
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 0
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 0
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 0
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 0
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_65
timestamp 0
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 0
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 0
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 0
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_97
timestamp 0
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_109
timestamp 0
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_121
timestamp 0
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_133
timestamp 0
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 0
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_141
timestamp 0
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_153
timestamp 0
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_165
timestamp 0
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_177
timestamp 0
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_189
timestamp 0
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 0
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 0
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_209
timestamp 0
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_221
timestamp 0
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_233
timestamp 0
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_245
timestamp 0
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_251
timestamp 0
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 0
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_265
timestamp 0
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_277
timestamp 0
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_289
timestamp 0
transform 1 0 27692 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_297
timestamp 0
transform 1 0 28428 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 0
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 0
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 0
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 0
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 0
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 0
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 0
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_69
timestamp 0
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_81
timestamp 0
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_93
timestamp 0
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_105
timestamp 0
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 0
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 0
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_125
timestamp 0
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_137
timestamp 0
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_149
timestamp 0
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_161
timestamp 0
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 0
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 0
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_181
timestamp 0
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_193
timestamp 0
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_205
timestamp 0
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_217
timestamp 0
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 0
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_225
timestamp 0
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_237
timestamp 0
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_249
timestamp 0
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_261
timestamp 0
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_273
timestamp 0
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 0
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 0
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_293
timestamp 0
transform 1 0 28060 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 0
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 0
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 0
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 0
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 0
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 0
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_65
timestamp 0
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 0
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 0
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 0
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_97
timestamp 0
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_109
timestamp 0
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_121
timestamp 0
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_133
timestamp 0
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 0
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_141
timestamp 0
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_153
timestamp 0
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_165
timestamp 0
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_177
timestamp 0
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_189
timestamp 0
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 0
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 0
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_209
timestamp 0
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_221
timestamp 0
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_233
timestamp 0
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_245
timestamp 0
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 0
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 0
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_265
timestamp 0
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_277
timestamp 0
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_289
timestamp 0
transform 1 0 27692 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_297
timestamp 0
transform 1 0 28428 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 0
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 0
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 0
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 0
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 0
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 0
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 0
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_69
timestamp 0
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_81
timestamp 0
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_93
timestamp 0
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_105
timestamp 0
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 0
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_113
timestamp 0
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_125
timestamp 0
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_137
timestamp 0
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_149
timestamp 0
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_161
timestamp 0
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 0
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 0
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_181
timestamp 0
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_193
timestamp 0
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_205
timestamp 0
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_217
timestamp 0
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 0
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 0
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_237
timestamp 0
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_249
timestamp 0
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_261
timestamp 0
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_273
timestamp 0
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 0
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 0
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_293
timestamp 0
transform 1 0 28060 0 -1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_3
timestamp 0
transform 1 0 1380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_15
timestamp 0
transform 1 0 2484 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 0
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 0
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 0
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 0
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 0
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 0
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 0
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 0
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_97
timestamp 0
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_109
timestamp 0
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_121
timestamp 0
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_133
timestamp 0
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 0
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_141
timestamp 0
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_153
timestamp 0
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_165
timestamp 0
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_177
timestamp 0
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_189
timestamp 0
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 0
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_197
timestamp 0
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_209
timestamp 0
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_221
timestamp 0
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_233
timestamp 0
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_245
timestamp 0
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 0
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 0
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_265
timestamp 0
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_277
timestamp 0
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 0
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 0
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 0
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 0
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 0
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 0
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 0
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 0
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_81
timestamp 0
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_93
timestamp 0
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_105
timestamp 0
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 0
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 0
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 0
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_137
timestamp 0
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_149
timestamp 0
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_161
timestamp 0
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 0
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 0
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_181
timestamp 0
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_193
timestamp 0
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_205
timestamp 0
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_217
timestamp 0
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_223
timestamp 0
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 0
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_237
timestamp 0
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_249
timestamp 0
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_261
timestamp 0
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_273
timestamp 0
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 0
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 0
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_293
timestamp 0
transform 1 0 28060 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 0
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 0
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 0
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 0
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 0
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 0
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 0
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 0
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 0
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 0
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 0
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_109
timestamp 0
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_121
timestamp 0
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_133
timestamp 0
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 0
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 0
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_153
timestamp 0
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_165
timestamp 0
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_177
timestamp 0
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_189
timestamp 0
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 0
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_197
timestamp 0
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_209
timestamp 0
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_221
timestamp 0
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_233
timestamp 0
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_245
timestamp 0
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 0
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 0
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 0
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_277
timestamp 0
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_289
timestamp 0
transform 1 0 27692 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_297
timestamp 0
transform 1 0 28428 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 0
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 0
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 0
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 0
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 0
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 0
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 0
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 0
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 0
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_93
timestamp 0
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 0
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 0
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 0
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_125
timestamp 0
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_137
timestamp 0
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_149
timestamp 0
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_161
timestamp 0
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 0
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 0
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_181
timestamp 0
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_193
timestamp 0
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_205
timestamp 0
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_217
timestamp 0
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 0
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 0
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_237
timestamp 0
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_249
timestamp 0
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_261
timestamp 0
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_273
timestamp 0
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_279
timestamp 0
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 0
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_293
timestamp 0
transform 1 0 28060 0 -1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_9
timestamp 0
transform 1 0 1932 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_21
timestamp 0
transform 1 0 3036 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 0
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 0
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 0
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_53
timestamp 0
transform 1 0 5980 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_57
timestamp 0
transform 1 0 6348 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_65
timestamp 0
transform 1 0 7084 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_72
timestamp 0
transform 1 0 7728 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 0
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 0
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_109
timestamp 0
transform 1 0 11132 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_113
timestamp 0
transform 1 0 11500 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_125
timestamp 0
transform 1 0 12604 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_137
timestamp 0
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 0
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_153
timestamp 0
transform 1 0 15180 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_161
timestamp 0
transform 1 0 15916 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_167
timestamp 0
transform 1 0 16468 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_169
timestamp 0
transform 1 0 16652 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_181
timestamp 0
transform 1 0 17756 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_193
timestamp 0
transform 1 0 18860 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 0
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_209
timestamp 0
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_221
timestamp 0
transform 1 0 21436 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_225
timestamp 0
transform 1 0 21804 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_237
timestamp 0
transform 1 0 22908 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_249
timestamp 0
transform 1 0 24012 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_253
timestamp 0
transform 1 0 24380 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_261
timestamp 0
transform 1 0 25116 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_272
timestamp 0
transform 1 0 26128 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_281
timestamp 0
transform 1 0 26956 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_293
timestamp 0
transform 1 0 28060 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 0
transform 1 0 19320 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 0
transform -1 0 25116 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 0
transform -1 0 25944 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 0
transform 1 0 21896 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 0
transform 1 0 21988 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 0
transform -1 0 23460 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 0
transform -1 0 25668 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 0
transform -1 0 19964 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 0
transform 1 0 18032 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 0
transform -1 0 24380 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 0
transform -1 0 21528 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 0
transform -1 0 19228 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 0
transform -1 0 18952 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 0
transform 1 0 17480 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 0
transform 1 0 17664 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 0
transform -1 0 19964 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 0
transform -1 0 16008 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 0
transform -1 0 26864 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 0
transform -1 0 19136 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 0
transform -1 0 18216 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 0
transform -1 0 16652 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 0
transform -1 0 18216 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 0
transform -1 0 18768 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 0
transform -1 0 20792 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 0
transform -1 0 16008 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 0
transform -1 0 16744 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 0
transform -1 0 18400 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input2
timestamp 0
transform 1 0 25208 0 1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input3
timestamp 0
transform 1 0 1380 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 0
transform -1 0 27416 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 0
transform 1 0 16192 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8
timestamp 0
transform -1 0 28612 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 0
transform 1 0 9108 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10
timestamp 0
transform -1 0 28612 0 -1 6528
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  output11
timestamp 0
transform -1 0 1932 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output12
timestamp 0
transform -1 0 7728 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 0
transform -1 0 28888 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 0
transform -1 0 28888 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 0
transform -1 0 28888 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 0
transform -1 0 28888 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 0
transform -1 0 28888 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 0
transform -1 0 28888 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 0
transform -1 0 28888 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 0
transform -1 0 28888 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 0
transform -1 0 28888 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 0
transform -1 0 28888 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 0
transform -1 0 28888 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 0
transform -1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 0
transform -1 0 28888 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 0
transform -1 0 28888 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 0
transform -1 0 28888 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 0
transform -1 0 28888 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 0
transform -1 0 28888 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 0
transform -1 0 28888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 0
transform -1 0 28888 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 0
transform -1 0 28888 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 0
transform -1 0 28888 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 0
transform -1 0 28888 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 0
transform -1 0 28888 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 0
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 0
transform -1 0 28888 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 0
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 0
transform -1 0 28888 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 0
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 0
transform -1 0 28888 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 0
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 0
transform -1 0 28888 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 0
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 0
transform -1 0 28888 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 0
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 0
transform -1 0 28888 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 0
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 0
transform -1 0 28888 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 0
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 0
transform -1 0 28888 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 0
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 0
transform -1 0 28888 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 0
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 0
transform -1 0 28888 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 0
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 0
transform -1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 0
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 0
transform -1 0 28888 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 0
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 0
transform -1 0 28888 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 0
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 0
transform -1 0 28888 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 0
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 0
transform -1 0 28888 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 0
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 0
transform -1 0 28888 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 0
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 0
transform -1 0 28888 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 0
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 0
transform -1 0 28888 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 0
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 0
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 0
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 0
transform -1 0 28888 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 0
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 0
transform -1 0 28888 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 0
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 0
transform -1 0 28888 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 0
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 0
transform -1 0 28888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 0
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 0
transform -1 0 28888 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 0
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 0
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 0
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 0
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 0
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 0
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 0
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 0
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 0
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 0
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 0
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 0
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 0
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 0
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 0
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 0
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 0
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 0
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 0
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 0
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 0
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 0
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 0
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 0
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 0
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 0
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 0
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 0
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 0
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 0
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 0
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 0
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 0
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 0
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 0
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 0
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 0
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 0
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 0
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 0
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 0
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 0
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 0
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 0
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 0
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 0
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 0
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 0
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 0
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 0
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 0
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 0
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 0
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 0
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 0
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 0
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 0
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 0
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 0
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 0
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 0
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 0
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 0
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 0
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 0
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 0
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 0
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 0
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 0
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 0
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 0
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 0
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 0
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 0
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 0
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 0
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 0
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 0
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 0
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 0
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 0
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 0
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 0
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 0
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 0
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 0
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 0
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 0
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 0
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 0
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 0
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 0
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 0
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 0
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 0
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 0
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 0
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 0
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 0
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 0
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 0
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 0
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 0
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 0
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 0
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 0
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 0
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 0
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 0
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 0
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 0
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 0
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 0
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 0
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 0
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 0
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 0
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 0
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 0
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 0
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 0
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 0
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 0
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 0
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 0
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 0
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 0
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 0
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 0
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 0
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 0
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 0
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 0
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 0
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 0
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 0
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 0
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 0
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 0
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 0
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 0
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 0
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 0
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 0
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 0
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 0
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 0
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 0
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 0
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 0
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 0
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 0
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 0
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 0
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 0
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 0
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 0
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 0
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 0
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 0
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 0
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 0
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 0
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 0
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 0
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 0
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 0
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 0
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 0
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 0
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 0
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 0
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 0
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 0
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 0
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 0
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 0
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 0
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 0
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 0
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 0
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 0
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 0
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 0
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 0
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 0
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 0
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 0
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 0
transform 1 0 6256 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 0
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 0
transform 1 0 11408 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 0
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 0
transform 1 0 16560 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 0
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 0
transform 1 0 21712 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 0
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 0
transform 1 0 26864 0 1 27200
box -38 -48 130 592
<< labels >>
rlabel metal1 s 14996 27200 14996 27200 4 VGND
rlabel metal1 s 14996 27744 14996 27744 4 VPWR
rlabel metal1 s 19228 10574 19228 10574 4 _000_
rlabel metal1 s 20286 9418 20286 9418 4 _001_
rlabel metal2 s 22494 10914 22494 10914 4 _002_
rlabel metal1 s 22862 10574 22862 10574 4 _003_
rlabel metal1 s 23598 8568 23598 8568 4 _004_
rlabel metal1 s 22770 9690 22770 9690 4 _005_
rlabel metal1 s 20148 2618 20148 2618 4 _006_
rlabel metal1 s 22080 2618 22080 2618 4 _007_
rlabel metal1 s 20976 4046 20976 4046 4 _008_
rlabel metal1 s 24610 3570 24610 3570 4 _009_
rlabel metal2 s 24702 4828 24702 4828 4 _010_
rlabel metal1 s 24472 5882 24472 5882 4 _011_
rlabel metal1 s 21252 5746 21252 5746 4 _012_
rlabel metal1 s 22457 6970 22457 6970 4 _013_
rlabel metal1 s 23552 6970 23552 6970 4 _014_
rlabel metal1 s 20010 6392 20010 6392 4 _015_
rlabel metal1 s 18170 3128 18170 3128 4 _016_
rlabel metal1 s 16238 4250 16238 4250 4 _017_
rlabel metal1 s 16974 5304 16974 5304 4 _018_
rlabel metal1 s 17066 3162 17066 3162 4 _019_
rlabel metal1 s 17618 4794 17618 4794 4 _020_
rlabel metal1 s 19504 4250 19504 4250 4 _021_
rlabel metal2 s 18722 7140 18722 7140 4 _022_
rlabel metal1 s 16875 6970 16875 6970 4 _023_
rlabel metal1 s 19918 8398 19918 8398 4 _024_
rlabel metal1 s 17756 10098 17756 10098 4 _025_
rlabel metal2 s 17342 10880 17342 10880 4 _026_
rlabel metal2 s 15042 10982 15042 10982 4 _027_
rlabel metal1 s 14674 9690 14674 9690 4 _028_
rlabel metal2 s 16238 8126 16238 8126 4 _029_
rlabel metal1 s 14168 8534 14168 8534 4 _030_
rlabel metal1 s 14812 11798 14812 11798 4 _031_
rlabel metal1 s 16146 12274 16146 12274 4 _032_
rlabel metal2 s 23690 4794 23690 4794 4 _033_
rlabel metal2 s 22770 6596 22770 6596 4 _034_
rlabel metal1 s 19826 5304 19826 5304 4 _035_
rlabel metal2 s 21942 6358 21942 6358 4 _036_
rlabel metal1 s 23046 2618 23046 2618 4 _037_
rlabel metal1 s 21252 7174 21252 7174 4 _038_
rlabel metal2 s 22494 8160 22494 8160 4 _039_
rlabel metal1 s 19826 9588 19826 9588 4 _040_
rlabel metal1 s 20930 8500 20930 8500 4 _041_
rlabel metal1 s 23276 8534 23276 8534 4 _042_
rlabel metal1 s 22770 9418 22770 9418 4 _043_
rlabel metal1 s 22264 9690 22264 9690 4 _044_
rlabel metal1 s 23046 2448 23046 2448 4 _045_
rlabel metal1 s 23368 8942 23368 8942 4 _046_
rlabel metal1 s 23598 8976 23598 8976 4 _047_
rlabel metal2 s 20738 7514 20738 7514 4 _048_
rlabel metal1 s 20516 3502 20516 3502 4 _049_
rlabel metal1 s 19596 2414 19596 2414 4 _050_
rlabel metal1 s 20608 2414 20608 2414 4 _051_
rlabel metal1 s 22218 2516 22218 2516 4 _052_
rlabel metal2 s 22678 2924 22678 2924 4 _053_
rlabel metal2 s 21942 4352 21942 4352 4 _054_
rlabel metal1 s 22034 4080 22034 4080 4 _055_
rlabel metal1 s 23460 3502 23460 3502 4 _056_
rlabel metal1 s 23092 5202 23092 5202 4 _057_
rlabel metal1 s 23690 3502 23690 3502 4 _058_
rlabel metal1 s 25438 5746 25438 5746 4 _059_
rlabel metal1 s 24564 5202 24564 5202 4 _060_
rlabel metal1 s 24610 5644 24610 5644 4 _061_
rlabel metal1 s 25116 5746 25116 5746 4 _062_
rlabel metal1 s 23414 5304 23414 5304 4 _063_
rlabel metal1 s 22218 5656 22218 5656 4 _064_
rlabel metal1 s 23782 6256 23782 6256 4 _065_
rlabel metal1 s 23782 6800 23782 6800 4 _066_
rlabel metal2 s 22678 6528 22678 6528 4 _067_
rlabel metal1 s 19826 5882 19826 5882 4 _068_
rlabel metal1 s 20516 2550 20516 2550 4 _069_
rlabel metal1 s 16836 4114 16836 4114 4 _070_
rlabel metal1 s 18400 3910 18400 3910 4 _071_
rlabel metal1 s 17434 3094 17434 3094 4 _072_
rlabel metal2 s 17986 5066 17986 5066 4 _073_
rlabel metal1 s 19642 4148 19642 4148 4 _074_
rlabel metal3 s 18722 7837 18722 7837 4 _075_
rlabel metal1 s 21068 7514 21068 7514 4 _076_
rlabel metal2 s 20562 8602 20562 8602 4 _077_
rlabel metal1 s 18400 6766 18400 6766 4 _078_
rlabel metal1 s 18078 7854 18078 7854 4 _079_
rlabel metal1 s 17664 7514 17664 7514 4 _080_
rlabel metal1 s 20746 8466 20746 8466 4 _081_
rlabel metal1 s 19780 8058 19780 8058 4 _082_
rlabel metal1 s 18492 10642 18492 10642 4 _083_
rlabel metal1 s 17388 10642 17388 10642 4 _084_
rlabel metal1 s 15088 10642 15088 10642 4 _085_
rlabel metal1 s 14996 9554 14996 9554 4 _086_
rlabel metal1 s 16376 8602 16376 8602 4 _087_
rlabel metal1 s 14352 8942 14352 8942 4 _088_
rlabel metal1 s 15318 12206 15318 12206 4 _089_
rlabel metal1 s 16698 12750 16698 12750 4 _090_
rlabel metal1 s 18722 12342 18722 12342 4 _091_
rlabel metal1 s 18814 12716 18814 12716 4 _092_
rlabel metal2 s 18952 11764 18952 11764 4 _093_
rlabel metal1 s 16146 9486 16146 9486 4 _094_
rlabel metal1 s 16698 10574 16698 10574 4 _095_
rlabel metal1 s 17756 10506 17756 10506 4 _096_
rlabel metal1 s 19504 11118 19504 11118 4 _097_
rlabel metal2 s 24150 8364 24150 8364 4 _098_
rlabel metal1 s 21436 8602 21436 8602 4 _099_
rlabel metal1 s 21298 8330 21298 8330 4 _100_
rlabel metal2 s 19274 11526 19274 11526 4 _101_
rlabel metal1 s 21390 9486 21390 9486 4 _102_
rlabel metal1 s 20102 8976 20102 8976 4 _103_
rlabel metal1 s 20378 9146 20378 9146 4 _104_
rlabel metal1 s 18814 9146 18814 9146 4 _105_
rlabel metal2 s 19642 9826 19642 9826 4 _106_
rlabel metal1 s 21206 9588 21206 9588 4 _107_
rlabel metal1 s 21528 9894 21528 9894 4 _108_
rlabel metal2 s 20562 9690 20562 9690 4 _109_
rlabel metal1 s 20884 9554 20884 9554 4 _110_
rlabel metal1 s 21206 9146 21206 9146 4 _111_
rlabel metal1 s 20056 7854 20056 7854 4 bit_idx\[0\]
rlabel metal2 s 19458 9248 19458 9248 4 bit_idx\[1\]
rlabel metal1 s 19366 8874 19366 8874 4 bit_idx\[2\]
rlabel metal3 s 24932 15640 24932 15640 4 clk
rlabel metal1 s 23184 2414 23184 2414 4 clk_cnt\[0\]
rlabel metal2 s 19918 4386 19918 4386 4 clk_cnt\[10\]
rlabel metal1 s 18216 4658 18216 4658 4 clk_cnt\[11\]
rlabel metal1 s 18768 5134 18768 5134 4 clk_cnt\[12\]
rlabel metal1 s 19182 4046 19182 4046 4 clk_cnt\[13\]
rlabel metal1 s 18906 6222 18906 6222 4 clk_cnt\[14\]
rlabel metal2 s 21022 5202 21022 5202 4 clk_cnt\[15\]
rlabel metal1 s 21574 4624 21574 4624 4 clk_cnt\[1\]
rlabel metal1 s 21758 4522 21758 4522 4 clk_cnt\[2\]
rlabel metal1 s 25898 4046 25898 4046 4 clk_cnt\[3\]
rlabel metal1 s 26036 5134 26036 5134 4 clk_cnt\[4\]
rlabel metal1 s 26358 6222 26358 6222 4 clk_cnt\[5\]
rlabel metal1 s 21942 5576 21942 5576 4 clk_cnt\[6\]
rlabel metal1 s 21942 6698 21942 6698 4 clk_cnt\[7\]
rlabel metal1 s 22954 7276 22954 7276 4 clk_cnt\[8\]
rlabel metal2 s 19826 5916 19826 5916 4 clk_cnt\[9\]
rlabel metal1 s 20700 8058 20700 8058 4 clknet_0_clk
rlabel metal1 s 17250 3570 17250 3570 4 clknet_2_0__leaf_clk
rlabel metal1 s 19918 11662 19918 11662 4 clknet_2_1__leaf_clk
rlabel metal2 s 21850 3196 21850 3196 4 clknet_2_2__leaf_clk
rlabel metal1 s 23322 7310 23322 7310 4 clknet_2_3__leaf_clk
rlabel metal2 s 18078 1588 18078 1588 4 data_in[0]
rlabel metal1 s 25208 27506 25208 27506 4 data_in[1]
rlabel metal3 s 820 18428 820 18428 4 data_in[2]
rlabel metal2 s 46 1588 46 1588 4 data_in[3]
rlabel metal2 s 27094 1588 27094 1588 4 data_in[4]
rlabel metal3 s 820 8908 820 8908 4 data_in[5]
rlabel metal1 s 16192 27438 16192 27438 4 data_in[6]
rlabel metal3 s 28566 25245 28566 25245 4 data_in[7]
rlabel metal1 s 18768 10098 18768 10098 4 data_reg\[0\]
rlabel metal1 s 18032 11254 18032 11254 4 data_reg\[1\]
rlabel metal1 s 16238 10574 16238 10574 4 data_reg\[2\]
rlabel metal2 s 17700 9486 17700 9486 4 data_reg\[3\]
rlabel metal1 s 16560 8942 16560 8942 4 data_reg\[4\]
rlabel metal1 s 16238 9010 16238 9010 4 data_reg\[5\]
rlabel metal1 s 16836 11594 16836 11594 4 data_reg\[6\]
rlabel metal1 s 17756 12750 17756 12750 4 data_reg\[7\]
rlabel metal1 s 17940 12274 17940 12274 4 net1
rlabel metal1 s 21942 8500 21942 8500 4 net10
rlabel metal1 s 4347 27370 4347 27370 4 net11
rlabel metal1 s 7498 27472 7498 27472 4 net12
rlabel metal2 s 19734 9078 19734 9078 4 net13
rlabel metal1 s 18591 9962 18591 9962 4 net14
rlabel metal1 s 21489 6698 21489 6698 4 net15
rlabel metal1 s 21114 2414 21114 2414 4 net16
rlabel metal1 s 20378 8534 20378 8534 4 net17
rlabel metal1 s 24196 6766 24196 6766 4 net18
rlabel metal1 s 24150 5236 24150 5236 4 net19
rlabel metal1 s 17710 12206 17710 12206 4 net2
rlabel metal1 s 22816 6766 22816 6766 4 net20
rlabel metal1 s 22586 4114 22586 4114 4 net21
rlabel metal1 s 22724 5678 22724 5678 4 net22
rlabel metal2 s 24978 4386 24978 4386 4 net23
rlabel metal1 s 18998 5746 18998 5746 4 net24
rlabel metal2 s 19366 4454 19366 4454 4 net25
rlabel metal1 s 22310 2380 22310 2380 4 net26
rlabel metal1 s 20792 5134 20792 5134 4 net27
rlabel metal1 s 17894 4046 17894 4046 4 net28
rlabel metal1 s 17618 4012 17618 4012 4 net29
rlabel metal1 s 7590 18734 7590 18734 4 net3
rlabel metal1 s 18400 5746 18400 5746 4 net30
rlabel metal2 s 18354 7752 18354 7752 4 net31
rlabel metal1 s 19320 3366 19320 3366 4 net32
rlabel metal1 s 15088 8806 15088 8806 4 net33
rlabel metal1 s 24702 5780 24702 5780 4 net34
rlabel metal1 s 18032 10778 18032 10778 4 net35
rlabel metal1 s 17342 8466 17342 8466 4 net36
rlabel metal1 s 14398 9588 14398 9588 4 net37
rlabel metal1 s 17342 12818 17342 12818 4 net38
rlabel metal1 s 17894 11730 17894 11730 4 net39
rlabel metal1 s 7636 2482 7636 2482 4 net4
rlabel metal1 s 19918 11050 19918 11050 4 net40
rlabel metal1 s 14904 10574 14904 10574 4 net41
rlabel metal1 s 16008 12954 16008 12954 4 net42
rlabel metal1 s 18032 2346 18032 2346 4 net5
rlabel metal1 s 4255 8806 4255 8806 4 net6
rlabel metal1 s 16974 12784 16974 12784 4 net7
rlabel metal1 s 18446 12852 18446 12852 4 net8
rlabel metal1 s 14076 2278 14076 2278 4 net9
rlabel metal1 s 20608 10778 20608 10778 4 parity_bit
rlabel metal2 s 9062 1027 9062 1027 4 rst_n
rlabel metal2 s 21114 9248 21114 9248 4 state\[0\]
rlabel metal1 s 24932 8330 24932 8330 4 state\[1\]
rlabel metal1 s 21804 9554 21804 9554 4 state\[2\]
rlabel metal3 s 0 27888 800 28008 4 tx_busy
port 13 nsew
rlabel metal1 s 7268 27574 7268 27574 4 tx_out
rlabel metal3 s 28566 6205 28566 6205 4 tx_start
flabel metal5 s 1056 25048 28936 25368 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 18656 28936 18976 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 12264 28936 12584 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 5872 28936 6192 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 25915 2128 26235 27792 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 18969 2128 19289 27792 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 12023 2128 12343 27792 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 5077 2128 5397 27792 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 1056 24388 28936 24708 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 17996 28936 18316 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 11604 28936 11924 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 5212 28936 5532 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 25255 2128 25575 27792 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 18309 2128 18629 27792 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 11363 2128 11683 27792 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 4417 2128 4737 27792 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 29200 15648 30000 15768 0 FreeSans 600 0 0 0 clk
port 3 nsew
flabel metal2 s 18050 0 18106 800 0 FreeSans 280 90 0 0 data_in[0]
port 4 nsew
flabel metal2 s 25134 29200 25190 30000 0 FreeSans 280 90 0 0 data_in[1]
port 5 nsew
flabel metal3 s 0 18368 800 18488 0 FreeSans 600 0 0 0 data_in[2]
port 6 nsew
flabel metal2 s 18 0 74 800 0 FreeSans 280 90 0 0 data_in[3]
port 7 nsew
flabel metal2 s 27066 0 27122 800 0 FreeSans 280 90 0 0 data_in[4]
port 8 nsew
flabel metal3 s 0 8848 800 8968 0 FreeSans 600 0 0 0 data_in[5]
port 9 nsew
flabel metal2 s 16118 29200 16174 30000 0 FreeSans 280 90 0 0 data_in[6]
port 10 nsew
flabel metal3 s 29200 25168 30000 25288 0 FreeSans 600 0 0 0 data_in[7]
port 11 nsew
flabel metal2 s 9034 0 9090 800 0 FreeSans 280 90 0 0 rst_n
port 12 nsew
flabel metal3 s 400 27948 400 27948 0 FreeSans 600 0 0 0 tx_busy
flabel metal2 s 7102 29200 7158 30000 0 FreeSans 280 90 0 0 tx_out
port 14 nsew
flabel metal3 s 29200 6128 30000 6248 0 FreeSans 600 0 0 0 tx_start
port 15 nsew
<< properties >>
string FIXED_BBOX 0 0 30000 30000
<< end >>
