magic
tech sky130A
magscale 1 2
timestamp 1765484971
<< checkpaint >>
rect -1260 -1260 41260 41260
<< viali >>
rect 1501 37417 1535 37451
rect 9873 37417 9907 37451
rect 22017 37281 22051 37315
rect 22293 37213 22327 37247
rect 33793 37213 33827 37247
rect 1777 37145 1811 37179
rect 10149 37145 10183 37179
rect 33701 37077 33735 37111
rect 38393 33473 38427 33507
rect 38301 33269 38335 33303
rect 1501 25177 1535 25211
rect 1685 25177 1719 25211
rect 23673 16065 23707 16099
rect 22845 15997 22879 16031
rect 23765 15997 23799 16031
rect 22293 15861 22327 15895
rect 23949 15861 23983 15895
rect 23765 15589 23799 15623
rect 22109 15521 22143 15555
rect 22201 15521 22235 15555
rect 23305 15521 23339 15555
rect 24501 15521 24535 15555
rect 20729 15453 20763 15487
rect 21373 15453 21407 15487
rect 23029 15453 23063 15487
rect 23397 15453 23431 15487
rect 24593 15453 24627 15487
rect 22017 15385 22051 15419
rect 20545 15317 20579 15351
rect 21189 15317 21223 15351
rect 21649 15317 21683 15351
rect 22477 15317 22511 15351
rect 24961 15317 24995 15351
rect 21833 15113 21867 15147
rect 22201 15113 22235 15147
rect 22293 15113 22327 15147
rect 23673 15113 23707 15147
rect 20177 15045 20211 15079
rect 18981 14977 19015 15011
rect 23121 14977 23155 15011
rect 23765 14977 23799 15011
rect 24133 14977 24167 15011
rect 25053 14977 25087 15011
rect 25697 14977 25731 15011
rect 19901 14909 19935 14943
rect 22385 14909 22419 14943
rect 23857 14909 23891 14943
rect 24777 14909 24811 14943
rect 24961 14909 24995 14943
rect 21649 14841 21683 14875
rect 23305 14841 23339 14875
rect 18797 14773 18831 14807
rect 22937 14773 22971 14807
rect 25329 14773 25363 14807
rect 25513 14773 25547 14807
rect 19257 14569 19291 14603
rect 22385 14569 22419 14603
rect 24225 14501 24259 14535
rect 19901 14433 19935 14467
rect 20637 14433 20671 14467
rect 22477 14433 22511 14467
rect 22753 14433 22787 14467
rect 25881 14433 25915 14467
rect 26157 14433 26191 14467
rect 28181 14433 28215 14467
rect 19625 14365 19659 14399
rect 25053 14365 25087 14399
rect 25697 14365 25731 14399
rect 20913 14297 20947 14331
rect 27905 14297 27939 14331
rect 19717 14229 19751 14263
rect 24409 14229 24443 14263
rect 25329 14229 25363 14263
rect 25789 14229 25823 14263
rect 20453 14025 20487 14059
rect 26985 14025 27019 14059
rect 27905 14025 27939 14059
rect 18889 13957 18923 13991
rect 25145 13957 25179 13991
rect 22017 13889 22051 13923
rect 22937 13889 22971 13923
rect 27721 13889 27755 13923
rect 18613 13821 18647 13855
rect 20361 13821 20395 13855
rect 21005 13821 21039 13855
rect 21925 13821 21959 13855
rect 23213 13821 23247 13855
rect 24869 13821 24903 13855
rect 26617 13821 26651 13855
rect 27537 13821 27571 13855
rect 22293 13685 22327 13719
rect 24685 13685 24719 13719
rect 19717 13481 19751 13515
rect 23213 13481 23247 13515
rect 27537 13481 27571 13515
rect 20821 13413 20855 13447
rect 23489 13413 23523 13447
rect 19533 13345 19567 13379
rect 20545 13345 20579 13379
rect 24041 13345 24075 13379
rect 24869 13345 24903 13379
rect 26985 13345 27019 13379
rect 27997 13345 28031 13379
rect 19441 13277 19475 13311
rect 20453 13277 20487 13311
rect 20913 13277 20947 13311
rect 23397 13277 23431 13311
rect 23857 13277 23891 13311
rect 23949 13277 23983 13311
rect 25237 13277 25271 13311
rect 27721 13277 27755 13311
rect 28089 13277 28123 13311
rect 21189 13209 21223 13243
rect 27169 13209 27203 13243
rect 22661 13141 22695 13175
rect 26663 13141 26697 13175
rect 27077 13141 27111 13175
rect 21281 12937 21315 12971
rect 19809 12869 19843 12903
rect 1409 12801 1443 12835
rect 19165 12801 19199 12835
rect 19901 12801 19935 12835
rect 20453 12801 20487 12835
rect 21465 12801 21499 12835
rect 22870 12801 22904 12835
rect 24409 12801 24443 12835
rect 25421 12801 25455 12835
rect 25697 12801 25731 12835
rect 25881 12801 25915 12835
rect 26065 12801 26099 12835
rect 26617 12801 26651 12835
rect 26801 12801 26835 12835
rect 20085 12733 20119 12767
rect 21097 12733 21131 12767
rect 21833 12733 21867 12767
rect 22017 12733 22051 12767
rect 22753 12733 22787 12767
rect 23029 12733 23063 12767
rect 24547 12733 24581 12767
rect 24685 12733 24719 12767
rect 25605 12733 25639 12767
rect 26249 12733 26283 12767
rect 27445 12733 27479 12767
rect 27721 12733 27755 12767
rect 29469 12733 29503 12767
rect 19441 12665 19475 12699
rect 22477 12665 22511 12699
rect 24961 12665 24995 12699
rect 26525 12665 26559 12699
rect 1593 12597 1627 12631
rect 19349 12597 19383 12631
rect 23673 12597 23707 12631
rect 23765 12597 23799 12631
rect 25789 12597 25823 12631
rect 21005 12393 21039 12427
rect 21557 12393 21591 12427
rect 24593 12393 24627 12427
rect 27997 12393 28031 12427
rect 18981 12257 19015 12291
rect 22109 12257 22143 12291
rect 22937 12257 22971 12291
rect 24225 12257 24259 12291
rect 25881 12257 25915 12291
rect 26157 12257 26191 12291
rect 26617 12257 26651 12291
rect 27445 12257 27479 12291
rect 18061 12189 18095 12223
rect 19257 12189 19291 12223
rect 21925 12189 21959 12223
rect 23857 12189 23891 12223
rect 24041 12189 24075 12223
rect 24501 12189 24535 12223
rect 25421 12189 25455 12223
rect 25605 12189 25639 12223
rect 26249 12189 26283 12223
rect 26893 12189 26927 12223
rect 27077 12189 27111 12223
rect 27261 12189 27295 12223
rect 27721 12189 27755 12223
rect 28181 12189 28215 12223
rect 19533 12121 19567 12155
rect 25513 12121 25547 12155
rect 25743 12121 25777 12155
rect 26525 12121 26559 12155
rect 18245 12053 18279 12087
rect 18337 12053 18371 12087
rect 18705 12053 18739 12087
rect 18797 12053 18831 12087
rect 22017 12053 22051 12087
rect 22385 12053 22419 12087
rect 24961 12053 24995 12087
rect 25237 12053 25271 12087
rect 25973 12053 26007 12087
rect 27629 12053 27663 12087
rect 20453 11849 20487 11883
rect 22293 11849 22327 11883
rect 26801 11849 26835 11883
rect 20545 11781 20579 11815
rect 20913 11781 20947 11815
rect 25881 11781 25915 11815
rect 26985 11781 27019 11815
rect 18705 11713 18739 11747
rect 22201 11713 22235 11747
rect 22661 11713 22695 11747
rect 22845 11713 22879 11747
rect 25605 11713 25639 11747
rect 26341 11713 26375 11747
rect 26433 11713 26467 11747
rect 27149 11711 27183 11745
rect 29653 11713 29687 11747
rect 18981 11645 19015 11679
rect 22477 11645 22511 11679
rect 23029 11645 23063 11679
rect 23305 11645 23339 11679
rect 25421 11645 25455 11679
rect 25881 11645 25915 11679
rect 26249 11645 26283 11679
rect 27353 11645 27387 11679
rect 27537 11645 27571 11679
rect 27813 11645 27847 11679
rect 29561 11645 29595 11679
rect 21833 11509 21867 11543
rect 22753 11509 22787 11543
rect 24777 11509 24811 11543
rect 24869 11509 24903 11543
rect 25697 11509 25731 11543
rect 29837 11509 29871 11543
rect 19625 11305 19659 11339
rect 25421 11305 25455 11339
rect 26249 11305 26283 11339
rect 27813 11305 27847 11339
rect 27905 11305 27939 11339
rect 29101 11305 29135 11339
rect 20269 11169 20303 11203
rect 20729 11169 20763 11203
rect 24133 11169 24167 11203
rect 25145 11169 25179 11203
rect 25605 11169 25639 11203
rect 25881 11169 25915 11203
rect 26525 11169 26559 11203
rect 27077 11169 27111 11203
rect 27169 11169 27203 11203
rect 29009 11169 29043 11203
rect 23029 11101 23063 11135
rect 23121 11101 23155 11135
rect 23489 11101 23523 11135
rect 23581 11101 23615 11135
rect 24685 11101 24719 11135
rect 24777 11101 24811 11135
rect 25053 11101 25087 11135
rect 25697 11101 25731 11135
rect 25789 11101 25823 11135
rect 26893 11101 26927 11135
rect 27537 11101 27571 11135
rect 27629 11101 27663 11135
rect 28089 11101 28123 11135
rect 28365 11101 28399 11135
rect 28549 11101 28583 11135
rect 28825 11101 28859 11135
rect 29101 11101 29135 11135
rect 29561 11101 29595 11135
rect 29653 11101 29687 11135
rect 29837 11101 29871 11135
rect 21005 11033 21039 11067
rect 22753 11033 22787 11067
rect 23213 11033 23247 11067
rect 23351 11033 23385 11067
rect 26065 11033 26099 11067
rect 26281 11033 26315 11067
rect 27261 11033 27295 11067
rect 22845 10965 22879 10999
rect 24409 10965 24443 10999
rect 24869 10965 24903 10999
rect 26433 10965 26467 10999
rect 26709 10965 26743 10999
rect 26801 10965 26835 10999
rect 28641 10965 28675 10999
rect 30021 10965 30055 10999
rect 21281 10761 21315 10795
rect 23581 10761 23615 10795
rect 23765 10761 23799 10795
rect 27353 10761 27387 10795
rect 27629 10761 27663 10795
rect 29561 10761 29595 10795
rect 22109 10693 22143 10727
rect 26249 10693 26283 10727
rect 27470 10693 27504 10727
rect 28089 10693 28123 10727
rect 21465 10625 21499 10659
rect 23949 10625 23983 10659
rect 24041 10625 24075 10659
rect 24317 10625 24351 10659
rect 26341 10625 26375 10659
rect 26985 10625 27019 10659
rect 21833 10557 21867 10591
rect 27261 10557 27295 10591
rect 27813 10557 27847 10591
rect 24225 10489 24259 10523
rect 24961 10421 24995 10455
rect 26525 10421 26559 10455
rect 21097 10217 21131 10251
rect 23489 10217 23523 10251
rect 27537 10217 27571 10251
rect 24501 10081 24535 10115
rect 24593 10081 24627 10115
rect 24777 10081 24811 10115
rect 25605 10081 25639 10115
rect 23305 10013 23339 10047
rect 23673 10013 23707 10047
rect 24685 10013 24719 10047
rect 25237 10013 25271 10047
rect 25329 10013 25363 10047
rect 25513 10013 25547 10047
rect 25697 10013 25731 10047
rect 25789 10013 25823 10047
rect 28089 10013 28123 10047
rect 28457 10013 28491 10047
rect 29561 10013 29595 10047
rect 30113 10013 30147 10047
rect 22569 9945 22603 9979
rect 23857 9945 23891 9979
rect 26065 9945 26099 9979
rect 28181 9945 28215 9979
rect 28273 9945 28307 9979
rect 28733 9945 28767 9979
rect 28917 9945 28951 9979
rect 22753 9877 22787 9911
rect 24961 9877 24995 9911
rect 25973 9877 26007 9911
rect 27905 9877 27939 9911
rect 28549 9877 28583 9911
rect 25697 9673 25731 9707
rect 25881 9673 25915 9707
rect 29193 9673 29227 9707
rect 25513 9605 25547 9639
rect 27721 9605 27755 9639
rect 25283 9571 25317 9605
rect 22293 9537 22327 9571
rect 22477 9537 22511 9571
rect 24869 9537 24903 9571
rect 25789 9537 25823 9571
rect 26065 9537 26099 9571
rect 26157 9537 26191 9571
rect 26249 9537 26283 9571
rect 26433 9537 26467 9571
rect 26525 9537 26559 9571
rect 26617 9537 26651 9571
rect 26801 9537 26835 9571
rect 26985 9537 27019 9571
rect 24317 9469 24351 9503
rect 24593 9469 24627 9503
rect 25053 9469 25087 9503
rect 27077 9469 27111 9503
rect 27445 9469 27479 9503
rect 27353 9401 27387 9435
rect 22109 9333 22143 9367
rect 22845 9333 22879 9367
rect 24685 9333 24719 9367
rect 25145 9333 25179 9367
rect 25329 9333 25363 9367
rect 26801 9333 26835 9367
rect 27169 9333 27203 9367
rect 22937 9129 22971 9163
rect 24133 9129 24167 9163
rect 28549 9129 28583 9163
rect 29837 9129 29871 9163
rect 23857 9061 23891 9095
rect 29561 9061 29595 9095
rect 21189 8993 21223 9027
rect 23213 8993 23247 9027
rect 26157 8993 26191 9027
rect 26893 8993 26927 9027
rect 27261 8993 27295 9027
rect 27629 8993 27663 9027
rect 28273 8993 28307 9027
rect 23949 8925 23983 8959
rect 26341 8925 26375 8959
rect 26985 8925 27019 8959
rect 27169 8925 27203 8959
rect 28365 8925 28399 8959
rect 28641 8925 28675 8959
rect 29837 8925 29871 8959
rect 30021 8925 30055 8959
rect 21465 8857 21499 8891
rect 25881 8857 25915 8891
rect 27721 8857 27755 8891
rect 27997 8857 28031 8891
rect 24409 8789 24443 8823
rect 27905 8789 27939 8823
rect 28089 8789 28123 8823
rect 28917 8789 28951 8823
rect 21465 8585 21499 8619
rect 25881 8585 25915 8619
rect 38301 8585 38335 8619
rect 26249 8517 26283 8551
rect 29653 8517 29687 8551
rect 30389 8517 30423 8551
rect 21649 8449 21683 8483
rect 21833 8449 21867 8483
rect 23857 8449 23891 8483
rect 24133 8449 24167 8483
rect 26157 8449 26191 8483
rect 26341 8449 26375 8483
rect 26459 8449 26493 8483
rect 27629 8449 27663 8483
rect 27721 8449 27755 8483
rect 27813 8449 27847 8483
rect 27997 8449 28031 8483
rect 29929 8449 29963 8483
rect 30205 8449 30239 8483
rect 30297 8449 30331 8483
rect 30573 8449 30607 8483
rect 38393 8449 38427 8483
rect 22109 8381 22143 8415
rect 24041 8381 24075 8415
rect 24409 8381 24443 8415
rect 25973 8381 26007 8415
rect 26617 8381 26651 8415
rect 26985 8381 27019 8415
rect 27721 8313 27755 8347
rect 23581 8245 23615 8279
rect 23673 8245 23707 8279
rect 28181 8245 28215 8279
rect 30021 8245 30055 8279
rect 21281 8041 21315 8075
rect 22661 8041 22695 8075
rect 23213 8041 23247 8075
rect 24133 8041 24167 8075
rect 27353 8041 27387 8075
rect 30205 8041 30239 8075
rect 30941 8041 30975 8075
rect 23121 7905 23155 7939
rect 23581 7905 23615 7939
rect 29561 7905 29595 7939
rect 22569 7837 22603 7871
rect 22845 7837 22879 7871
rect 23213 7837 23247 7871
rect 25973 7837 26007 7871
rect 26065 7837 26099 7871
rect 27997 7837 28031 7871
rect 28089 7837 28123 7871
rect 28365 7837 28399 7871
rect 29009 7837 29043 7871
rect 29929 7837 29963 7871
rect 30021 7837 30055 7871
rect 30297 7837 30331 7871
rect 22937 7769 22971 7803
rect 23397 7701 23431 7735
rect 25789 7701 25823 7735
rect 28273 7701 28307 7735
rect 24041 7497 24075 7531
rect 26985 7497 27019 7531
rect 28365 7497 28399 7531
rect 30297 7497 30331 7531
rect 21281 7429 21315 7463
rect 20729 7361 20763 7395
rect 21005 7361 21039 7395
rect 21465 7361 21499 7395
rect 22017 7361 22051 7395
rect 23581 7361 23615 7395
rect 23857 7361 23891 7395
rect 24317 7361 24351 7395
rect 24409 7361 24443 7395
rect 24777 7361 24811 7395
rect 26525 7361 26559 7395
rect 26617 7361 26651 7395
rect 26801 7361 26835 7395
rect 27261 7361 27295 7395
rect 27445 7361 27479 7395
rect 28273 7361 28307 7395
rect 28457 7361 28491 7395
rect 28549 7361 28583 7395
rect 20821 7293 20855 7327
rect 21189 7293 21223 7327
rect 21649 7293 21683 7327
rect 22109 7293 22143 7327
rect 22753 7293 22787 7327
rect 23489 7293 23523 7327
rect 23673 7293 23707 7327
rect 27169 7293 27203 7327
rect 27353 7293 27387 7327
rect 27813 7293 27847 7327
rect 27905 7293 27939 7327
rect 27997 7293 28031 7327
rect 28089 7293 28123 7327
rect 28825 7293 28859 7327
rect 22845 7225 22879 7259
rect 27629 7225 27663 7259
rect 20545 7157 20579 7191
rect 21833 7157 21867 7191
rect 23581 7157 23615 7191
rect 24133 7157 24167 7191
rect 24593 7157 24627 7191
rect 26709 7157 26743 7191
rect 20440 6953 20474 6987
rect 24869 6953 24903 6987
rect 26985 6953 27019 6987
rect 27905 6953 27939 6987
rect 28641 6953 28675 6987
rect 29561 6953 29595 6987
rect 29837 6953 29871 6987
rect 29009 6885 29043 6919
rect 20177 6817 20211 6851
rect 21925 6817 21959 6851
rect 23673 6817 23707 6851
rect 24225 6817 24259 6851
rect 24777 6817 24811 6851
rect 25421 6817 25455 6851
rect 22477 6749 22511 6783
rect 22661 6749 22695 6783
rect 23305 6749 23339 6783
rect 24593 6749 24627 6783
rect 25329 6749 25363 6783
rect 25881 6749 25915 6783
rect 26065 6749 26099 6783
rect 26203 6749 26237 6783
rect 26341 6749 26375 6783
rect 26433 6749 26467 6783
rect 26617 6749 26651 6783
rect 26893 6749 26927 6783
rect 27261 6749 27295 6783
rect 27353 6749 27387 6783
rect 27813 6749 27847 6783
rect 28332 6749 28366 6783
rect 28733 6749 28767 6783
rect 28825 6749 28859 6783
rect 29837 6749 29871 6783
rect 30021 6749 30055 6783
rect 22109 6681 22143 6715
rect 23213 6681 23247 6715
rect 25237 6681 25271 6715
rect 25973 6681 26007 6715
rect 26801 6681 26835 6715
rect 27537 6681 27571 6715
rect 28549 6681 28583 6715
rect 23489 6613 23523 6647
rect 24409 6613 24443 6647
rect 25697 6613 25731 6647
rect 27169 6613 27203 6647
rect 28273 6613 28307 6647
rect 28457 6613 28491 6647
rect 21649 6409 21683 6443
rect 23673 6409 23707 6443
rect 25513 6409 25547 6443
rect 25881 6409 25915 6443
rect 26985 6409 27019 6443
rect 27721 6409 27755 6443
rect 24041 6341 24075 6375
rect 19901 6273 19935 6307
rect 25789 6273 25823 6307
rect 26801 6273 26835 6307
rect 29469 6273 29503 6307
rect 20177 6205 20211 6239
rect 21925 6205 21959 6239
rect 22201 6205 22235 6239
rect 23765 6205 23799 6239
rect 26525 6205 26559 6239
rect 27537 6205 27571 6239
rect 29193 6205 29227 6239
rect 26249 6069 26283 6103
rect 26525 6069 26559 6103
rect 22201 5865 22235 5899
rect 26157 5865 26191 5899
rect 27997 5865 28031 5899
rect 28917 5865 28951 5899
rect 23673 5729 23707 5763
rect 23949 5729 23983 5763
rect 24409 5729 24443 5763
rect 24685 5729 24719 5763
rect 26249 5729 26283 5763
rect 28825 5661 28859 5695
rect 28917 5661 28951 5695
rect 29193 5661 29227 5695
rect 26525 5593 26559 5627
rect 28181 5525 28215 5559
rect 29101 5525 29135 5559
rect 22477 5321 22511 5355
rect 25973 5321 26007 5355
rect 26617 5321 26651 5355
rect 28549 5321 28583 5355
rect 22661 5185 22695 5219
rect 26341 5185 26375 5219
rect 27169 5185 27203 5219
rect 27813 5185 27847 5219
rect 28457 5185 28491 5219
rect 26433 5117 26467 5151
rect 27261 4777 27295 4811
rect 26985 4709 27019 4743
rect 27261 4573 27295 4607
rect 27445 4573 27479 4607
rect 23949 2601 23983 2635
rect 24133 2397 24167 2431
rect 1501 2329 1535 2363
rect 1685 2329 1719 2363
rect 11805 2329 11839 2363
rect 11989 2329 12023 2363
rect 35541 2329 35575 2363
rect 35725 2329 35759 2363
<< metal1 >>
rect 1104 37562 38824 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38824 37562
rect 1104 37488 38824 37510
rect 934 37408 940 37460
rect 992 37448 998 37460
rect 1489 37451 1547 37457
rect 1489 37448 1501 37451
rect 992 37420 1501 37448
rect 992 37408 998 37420
rect 1489 37417 1501 37420
rect 1535 37417 1547 37451
rect 1489 37411 1547 37417
rect 9674 37408 9680 37460
rect 9732 37448 9738 37460
rect 9861 37451 9919 37457
rect 9861 37448 9873 37451
rect 9732 37420 9873 37448
rect 9732 37408 9738 37420
rect 9861 37417 9873 37420
rect 9907 37417 9919 37451
rect 9861 37411 9919 37417
rect 21910 37272 21916 37324
rect 21968 37312 21974 37324
rect 22005 37315 22063 37321
rect 22005 37312 22017 37315
rect 21968 37284 22017 37312
rect 21968 37272 21974 37284
rect 22005 37281 22017 37284
rect 22051 37281 22063 37315
rect 22005 37275 22063 37281
rect 22278 37204 22284 37256
rect 22336 37204 22342 37256
rect 33502 37204 33508 37256
rect 33560 37244 33566 37256
rect 33781 37247 33839 37253
rect 33781 37244 33793 37247
rect 33560 37216 33793 37244
rect 33560 37204 33566 37216
rect 33781 37213 33793 37216
rect 33827 37213 33839 37247
rect 33781 37207 33839 37213
rect 1765 37179 1823 37185
rect 1765 37145 1777 37179
rect 1811 37176 1823 37179
rect 1811 37148 6914 37176
rect 1811 37145 1823 37148
rect 1765 37139 1823 37145
rect 6886 37108 6914 37148
rect 10134 37136 10140 37188
rect 10192 37136 10198 37188
rect 26234 37176 26240 37188
rect 16546 37148 26240 37176
rect 16546 37108 16574 37148
rect 26234 37136 26240 37148
rect 26292 37136 26298 37188
rect 6886 37080 16574 37108
rect 33686 37068 33692 37120
rect 33744 37068 33750 37120
rect 1104 37018 38824 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 35594 37018
rect 35646 36966 35658 37018
rect 35710 36966 35722 37018
rect 35774 36966 35786 37018
rect 35838 36966 35850 37018
rect 35902 36966 38824 37018
rect 1104 36944 38824 36966
rect 1104 36474 38824 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38824 36474
rect 1104 36400 38824 36422
rect 1104 35930 38824 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 35594 35930
rect 35646 35878 35658 35930
rect 35710 35878 35722 35930
rect 35774 35878 35786 35930
rect 35838 35878 35850 35930
rect 35902 35878 38824 35930
rect 1104 35856 38824 35878
rect 1104 35386 38824 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38824 35386
rect 1104 35312 38824 35334
rect 1104 34842 38824 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 35594 34842
rect 35646 34790 35658 34842
rect 35710 34790 35722 34842
rect 35774 34790 35786 34842
rect 35838 34790 35850 34842
rect 35902 34790 38824 34842
rect 1104 34768 38824 34790
rect 1104 34298 38824 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38824 34298
rect 1104 34224 38824 34246
rect 1104 33754 38824 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 35594 33754
rect 35646 33702 35658 33754
rect 35710 33702 35722 33754
rect 35774 33702 35786 33754
rect 35838 33702 35850 33754
rect 35902 33702 38824 33754
rect 1104 33680 38824 33702
rect 38381 33507 38439 33513
rect 38381 33473 38393 33507
rect 38427 33504 38439 33507
rect 38838 33504 38844 33516
rect 38427 33476 38844 33504
rect 38427 33473 38439 33476
rect 38381 33467 38439 33473
rect 38838 33464 38844 33476
rect 38896 33464 38902 33516
rect 38286 33260 38292 33312
rect 38344 33260 38350 33312
rect 1104 33210 38824 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38824 33210
rect 1104 33136 38824 33158
rect 1104 32666 38824 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 35594 32666
rect 35646 32614 35658 32666
rect 35710 32614 35722 32666
rect 35774 32614 35786 32666
rect 35838 32614 35850 32666
rect 35902 32614 38824 32666
rect 1104 32592 38824 32614
rect 1104 32122 38824 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38824 32122
rect 1104 32048 38824 32070
rect 1104 31578 38824 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 35594 31578
rect 35646 31526 35658 31578
rect 35710 31526 35722 31578
rect 35774 31526 35786 31578
rect 35838 31526 35850 31578
rect 35902 31526 38824 31578
rect 1104 31504 38824 31526
rect 1104 31034 38824 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38824 31034
rect 1104 30960 38824 30982
rect 1104 30490 38824 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 35594 30490
rect 35646 30438 35658 30490
rect 35710 30438 35722 30490
rect 35774 30438 35786 30490
rect 35838 30438 35850 30490
rect 35902 30438 38824 30490
rect 1104 30416 38824 30438
rect 1104 29946 38824 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38824 29946
rect 1104 29872 38824 29894
rect 1104 29402 38824 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 35594 29402
rect 35646 29350 35658 29402
rect 35710 29350 35722 29402
rect 35774 29350 35786 29402
rect 35838 29350 35850 29402
rect 35902 29350 38824 29402
rect 1104 29328 38824 29350
rect 1104 28858 38824 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38824 28858
rect 1104 28784 38824 28806
rect 1104 28314 38824 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 35594 28314
rect 35646 28262 35658 28314
rect 35710 28262 35722 28314
rect 35774 28262 35786 28314
rect 35838 28262 35850 28314
rect 35902 28262 38824 28314
rect 1104 28240 38824 28262
rect 1104 27770 38824 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38824 27770
rect 1104 27696 38824 27718
rect 1104 27226 38824 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 35594 27226
rect 35646 27174 35658 27226
rect 35710 27174 35722 27226
rect 35774 27174 35786 27226
rect 35838 27174 35850 27226
rect 35902 27174 38824 27226
rect 1104 27152 38824 27174
rect 1104 26682 38824 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38824 26682
rect 1104 26608 38824 26630
rect 1104 26138 38824 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 35594 26138
rect 35646 26086 35658 26138
rect 35710 26086 35722 26138
rect 35774 26086 35786 26138
rect 35838 26086 35850 26138
rect 35902 26086 38824 26138
rect 1104 26064 38824 26086
rect 1104 25594 38824 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38824 25594
rect 1104 25520 38824 25542
rect 934 25168 940 25220
rect 992 25208 998 25220
rect 1489 25211 1547 25217
rect 1489 25208 1501 25211
rect 992 25180 1501 25208
rect 992 25168 998 25180
rect 1489 25177 1501 25180
rect 1535 25177 1547 25211
rect 1489 25171 1547 25177
rect 1673 25211 1731 25217
rect 1673 25177 1685 25211
rect 1719 25208 1731 25211
rect 1719 25180 6914 25208
rect 1719 25177 1731 25180
rect 1673 25171 1731 25177
rect 6886 25140 6914 25180
rect 19610 25140 19616 25152
rect 6886 25112 19616 25140
rect 19610 25100 19616 25112
rect 19668 25100 19674 25152
rect 1104 25050 38824 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 35594 25050
rect 35646 24998 35658 25050
rect 35710 24998 35722 25050
rect 35774 24998 35786 25050
rect 35838 24998 35850 25050
rect 35902 24998 38824 25050
rect 1104 24976 38824 24998
rect 1104 24506 38824 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38824 24506
rect 1104 24432 38824 24454
rect 1104 23962 38824 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 35594 23962
rect 35646 23910 35658 23962
rect 35710 23910 35722 23962
rect 35774 23910 35786 23962
rect 35838 23910 35850 23962
rect 35902 23910 38824 23962
rect 1104 23888 38824 23910
rect 1104 23418 38824 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38824 23418
rect 1104 23344 38824 23366
rect 1104 22874 38824 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 35594 22874
rect 35646 22822 35658 22874
rect 35710 22822 35722 22874
rect 35774 22822 35786 22874
rect 35838 22822 35850 22874
rect 35902 22822 38824 22874
rect 1104 22800 38824 22822
rect 1104 22330 38824 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38824 22330
rect 1104 22256 38824 22278
rect 1104 21786 38824 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 35594 21786
rect 35646 21734 35658 21786
rect 35710 21734 35722 21786
rect 35774 21734 35786 21786
rect 35838 21734 35850 21786
rect 35902 21734 38824 21786
rect 1104 21712 38824 21734
rect 1104 21242 38824 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38824 21242
rect 1104 21168 38824 21190
rect 1104 20698 38824 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 35594 20698
rect 35646 20646 35658 20698
rect 35710 20646 35722 20698
rect 35774 20646 35786 20698
rect 35838 20646 35850 20698
rect 35902 20646 38824 20698
rect 1104 20624 38824 20646
rect 1104 20154 38824 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38824 20154
rect 1104 20080 38824 20102
rect 1104 19610 38824 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 35594 19610
rect 35646 19558 35658 19610
rect 35710 19558 35722 19610
rect 35774 19558 35786 19610
rect 35838 19558 35850 19610
rect 35902 19558 38824 19610
rect 1104 19536 38824 19558
rect 1104 19066 38824 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38824 19066
rect 1104 18992 38824 19014
rect 1104 18522 38824 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 35594 18522
rect 35646 18470 35658 18522
rect 35710 18470 35722 18522
rect 35774 18470 35786 18522
rect 35838 18470 35850 18522
rect 35902 18470 38824 18522
rect 1104 18448 38824 18470
rect 1104 17978 38824 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38824 17978
rect 1104 17904 38824 17926
rect 1104 17434 38824 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 35594 17434
rect 35646 17382 35658 17434
rect 35710 17382 35722 17434
rect 35774 17382 35786 17434
rect 35838 17382 35850 17434
rect 35902 17382 38824 17434
rect 1104 17360 38824 17382
rect 1104 16890 38824 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38824 16890
rect 1104 16816 38824 16838
rect 1104 16346 38824 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 35594 16346
rect 35646 16294 35658 16346
rect 35710 16294 35722 16346
rect 35774 16294 35786 16346
rect 35838 16294 35850 16346
rect 35902 16294 38824 16346
rect 1104 16272 38824 16294
rect 23658 16056 23664 16108
rect 23716 16096 23722 16108
rect 33686 16096 33692 16108
rect 23716 16068 33692 16096
rect 23716 16056 23722 16068
rect 33686 16056 33692 16068
rect 33744 16056 33750 16108
rect 22370 15988 22376 16040
rect 22428 16028 22434 16040
rect 22833 16031 22891 16037
rect 22833 16028 22845 16031
rect 22428 16000 22845 16028
rect 22428 15988 22434 16000
rect 22833 15997 22845 16000
rect 22879 15997 22891 16031
rect 22833 15991 22891 15997
rect 23753 16031 23811 16037
rect 23753 15997 23765 16031
rect 23799 16028 23811 16031
rect 24210 16028 24216 16040
rect 23799 16000 24216 16028
rect 23799 15997 23811 16000
rect 23753 15991 23811 15997
rect 24210 15988 24216 16000
rect 24268 15988 24274 16040
rect 22278 15852 22284 15904
rect 22336 15852 22342 15904
rect 23934 15852 23940 15904
rect 23992 15852 23998 15904
rect 1104 15802 38824 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38824 15802
rect 1104 15728 38824 15750
rect 22278 15648 22284 15700
rect 22336 15648 22342 15700
rect 23934 15648 23940 15700
rect 23992 15648 23998 15700
rect 22296 15620 22324 15648
rect 22112 15592 22324 15620
rect 23753 15623 23811 15629
rect 22112 15561 22140 15592
rect 23753 15589 23765 15623
rect 23799 15589 23811 15623
rect 23952 15620 23980 15648
rect 23952 15592 24624 15620
rect 23753 15583 23811 15589
rect 22097 15555 22155 15561
rect 22097 15521 22109 15555
rect 22143 15521 22155 15555
rect 22097 15515 22155 15521
rect 22189 15555 22247 15561
rect 22189 15521 22201 15555
rect 22235 15521 22247 15555
rect 22189 15515 22247 15521
rect 20717 15487 20775 15493
rect 20717 15453 20729 15487
rect 20763 15484 20775 15487
rect 21082 15484 21088 15496
rect 20763 15456 21088 15484
rect 20763 15453 20775 15456
rect 20717 15447 20775 15453
rect 21082 15444 21088 15456
rect 21140 15444 21146 15496
rect 21361 15487 21419 15493
rect 21361 15453 21373 15487
rect 21407 15484 21419 15487
rect 21407 15456 21680 15484
rect 21407 15453 21419 15456
rect 21361 15447 21419 15453
rect 20530 15308 20536 15360
rect 20588 15308 20594 15360
rect 21174 15308 21180 15360
rect 21232 15308 21238 15360
rect 21652 15357 21680 15456
rect 21910 15444 21916 15496
rect 21968 15484 21974 15496
rect 22204 15484 22232 15515
rect 22278 15512 22284 15564
rect 22336 15552 22342 15564
rect 23293 15555 23351 15561
rect 23293 15552 23305 15555
rect 22336 15524 23305 15552
rect 22336 15512 22342 15524
rect 23293 15521 23305 15524
rect 23339 15521 23351 15555
rect 23768 15552 23796 15583
rect 24489 15555 24547 15561
rect 24489 15552 24501 15555
rect 23768 15524 24501 15552
rect 23293 15515 23351 15521
rect 24489 15521 24501 15524
rect 24535 15521 24547 15555
rect 24489 15515 24547 15521
rect 21968 15456 22232 15484
rect 21968 15444 21974 15456
rect 22922 15444 22928 15496
rect 22980 15484 22986 15496
rect 24596 15493 24624 15592
rect 23017 15487 23075 15493
rect 23017 15484 23029 15487
rect 22980 15456 23029 15484
rect 22980 15444 22986 15456
rect 23017 15453 23029 15456
rect 23063 15453 23075 15487
rect 23017 15447 23075 15453
rect 23385 15487 23443 15493
rect 23385 15453 23397 15487
rect 23431 15453 23443 15487
rect 23385 15447 23443 15453
rect 24581 15487 24639 15493
rect 24581 15453 24593 15487
rect 24627 15453 24639 15487
rect 38286 15484 38292 15496
rect 24581 15447 24639 15453
rect 26206 15456 38292 15484
rect 22005 15419 22063 15425
rect 22005 15385 22017 15419
rect 22051 15416 22063 15419
rect 23400 15416 23428 15447
rect 26206 15416 26234 15456
rect 38286 15444 38292 15456
rect 38344 15444 38350 15496
rect 22051 15388 26234 15416
rect 22051 15385 22063 15388
rect 22005 15379 22063 15385
rect 21637 15351 21695 15357
rect 21637 15317 21649 15351
rect 21683 15317 21695 15351
rect 21637 15311 21695 15317
rect 22462 15308 22468 15360
rect 22520 15308 22526 15360
rect 24946 15308 24952 15360
rect 25004 15308 25010 15360
rect 1104 15258 38824 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 35594 15258
rect 35646 15206 35658 15258
rect 35710 15206 35722 15258
rect 35774 15206 35786 15258
rect 35838 15206 35850 15258
rect 35902 15206 38824 15258
rect 1104 15184 38824 15206
rect 20530 15104 20536 15156
rect 20588 15104 20594 15156
rect 21082 15104 21088 15156
rect 21140 15144 21146 15156
rect 21821 15147 21879 15153
rect 21821 15144 21833 15147
rect 21140 15116 21833 15144
rect 21140 15104 21146 15116
rect 21821 15113 21833 15116
rect 21867 15113 21879 15147
rect 21821 15107 21879 15113
rect 22186 15104 22192 15156
rect 22244 15104 22250 15156
rect 22281 15147 22339 15153
rect 22281 15113 22293 15147
rect 22327 15144 22339 15147
rect 22462 15144 22468 15156
rect 22327 15116 22468 15144
rect 22327 15113 22339 15116
rect 22281 15107 22339 15113
rect 22462 15104 22468 15116
rect 22520 15104 22526 15156
rect 23658 15104 23664 15156
rect 23716 15104 23722 15156
rect 24946 15104 24952 15156
rect 25004 15104 25010 15156
rect 20165 15079 20223 15085
rect 20165 15045 20177 15079
rect 20211 15076 20223 15079
rect 20548 15076 20576 15104
rect 20211 15048 20576 15076
rect 22388 15048 23428 15076
rect 20211 15045 20223 15048
rect 20165 15039 20223 15045
rect 18966 14968 18972 15020
rect 19024 14968 19030 15020
rect 22278 15008 22284 15020
rect 21298 14980 22284 15008
rect 22278 14968 22284 14980
rect 22336 14968 22342 15020
rect 19889 14943 19947 14949
rect 19889 14909 19901 14943
rect 19935 14909 19947 14943
rect 19889 14903 19947 14909
rect 18782 14764 18788 14816
rect 18840 14764 18846 14816
rect 19904 14804 19932 14903
rect 20530 14900 20536 14952
rect 20588 14940 20594 14952
rect 21910 14940 21916 14952
rect 20588 14912 21916 14940
rect 20588 14900 20594 14912
rect 21910 14900 21916 14912
rect 21968 14940 21974 14952
rect 22388 14949 22416 15048
rect 23109 15011 23167 15017
rect 23109 14977 23121 15011
rect 23155 15008 23167 15011
rect 23155 14980 23336 15008
rect 23155 14977 23167 14980
rect 23109 14971 23167 14977
rect 22373 14943 22431 14949
rect 22373 14940 22385 14943
rect 21968 14912 22385 14940
rect 21968 14900 21974 14912
rect 22373 14909 22385 14912
rect 22419 14909 22431 14943
rect 22373 14903 22431 14909
rect 22922 14900 22928 14952
rect 22980 14900 22986 14952
rect 21637 14875 21695 14881
rect 21637 14841 21649 14875
rect 21683 14872 21695 14875
rect 22940 14872 22968 14900
rect 23308 14881 23336 14980
rect 23400 14940 23428 15048
rect 23753 15011 23811 15017
rect 23753 14977 23765 15011
rect 23799 15008 23811 15011
rect 24121 15011 24179 15017
rect 24121 15008 24133 15011
rect 23799 14980 24133 15008
rect 23799 14977 23811 14980
rect 23753 14971 23811 14977
rect 24121 14977 24133 14980
rect 24167 14977 24179 15011
rect 24121 14971 24179 14977
rect 24486 14968 24492 15020
rect 24544 15008 24550 15020
rect 24964 15008 24992 15104
rect 25041 15011 25099 15017
rect 25041 15008 25053 15011
rect 24544 14980 24900 15008
rect 24964 14980 25053 15008
rect 24544 14968 24550 14980
rect 23845 14943 23903 14949
rect 23845 14940 23857 14943
rect 23400 14912 23857 14940
rect 23845 14909 23857 14912
rect 23891 14940 23903 14943
rect 24026 14940 24032 14952
rect 23891 14912 24032 14940
rect 23891 14909 23903 14912
rect 23845 14903 23903 14909
rect 24026 14900 24032 14912
rect 24084 14900 24090 14952
rect 24765 14943 24823 14949
rect 24765 14909 24777 14943
rect 24811 14909 24823 14943
rect 24872 14940 24900 14980
rect 25041 14977 25053 14980
rect 25087 14977 25099 15011
rect 25041 14971 25099 14977
rect 25406 14968 25412 15020
rect 25464 15008 25470 15020
rect 25685 15011 25743 15017
rect 25685 15008 25697 15011
rect 25464 14980 25697 15008
rect 25464 14968 25470 14980
rect 25685 14977 25697 14980
rect 25731 14977 25743 15011
rect 25685 14971 25743 14977
rect 24949 14943 25007 14949
rect 24949 14940 24961 14943
rect 24872 14912 24961 14940
rect 24765 14903 24823 14909
rect 24949 14909 24961 14912
rect 24995 14909 25007 14943
rect 24949 14903 25007 14909
rect 21683 14844 22968 14872
rect 23293 14875 23351 14881
rect 21683 14841 21695 14844
rect 21637 14835 21695 14841
rect 23293 14841 23305 14875
rect 23339 14841 23351 14875
rect 24780 14872 24808 14903
rect 24780 14844 25084 14872
rect 23293 14835 23351 14841
rect 25056 14816 25084 14844
rect 20714 14804 20720 14816
rect 19904 14776 20720 14804
rect 20714 14764 20720 14776
rect 20772 14764 20778 14816
rect 22830 14764 22836 14816
rect 22888 14804 22894 14816
rect 22925 14807 22983 14813
rect 22925 14804 22937 14807
rect 22888 14776 22937 14804
rect 22888 14764 22894 14776
rect 22925 14773 22937 14776
rect 22971 14773 22983 14807
rect 22925 14767 22983 14773
rect 25038 14764 25044 14816
rect 25096 14764 25102 14816
rect 25314 14764 25320 14816
rect 25372 14764 25378 14816
rect 25498 14764 25504 14816
rect 25556 14764 25562 14816
rect 1104 14714 38824 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38824 14714
rect 1104 14640 38824 14662
rect 18966 14560 18972 14612
rect 19024 14600 19030 14612
rect 19245 14603 19303 14609
rect 19245 14600 19257 14603
rect 19024 14572 19257 14600
rect 19024 14560 19030 14572
rect 19245 14569 19257 14572
rect 19291 14569 19303 14603
rect 19245 14563 19303 14569
rect 20714 14560 20720 14612
rect 20772 14560 20778 14612
rect 22370 14560 22376 14612
rect 22428 14560 22434 14612
rect 19889 14467 19947 14473
rect 19889 14433 19901 14467
rect 19935 14464 19947 14467
rect 20070 14464 20076 14476
rect 19935 14436 20076 14464
rect 19935 14433 19947 14436
rect 19889 14427 19947 14433
rect 20070 14424 20076 14436
rect 20128 14464 20134 14476
rect 20530 14464 20536 14476
rect 20128 14436 20536 14464
rect 20128 14424 20134 14436
rect 20530 14424 20536 14436
rect 20588 14424 20594 14476
rect 20625 14467 20683 14473
rect 20625 14433 20637 14467
rect 20671 14464 20683 14467
rect 20732 14464 20760 14560
rect 24213 14535 24271 14541
rect 24213 14501 24225 14535
rect 24259 14532 24271 14535
rect 25038 14532 25044 14544
rect 24259 14504 25044 14532
rect 24259 14501 24271 14504
rect 24213 14495 24271 14501
rect 25038 14492 25044 14504
rect 25096 14492 25102 14544
rect 21910 14464 21916 14476
rect 20671 14436 21916 14464
rect 20671 14433 20683 14436
rect 20625 14427 20683 14433
rect 21910 14424 21916 14436
rect 21968 14464 21974 14476
rect 22465 14467 22523 14473
rect 22465 14464 22477 14467
rect 21968 14436 22477 14464
rect 21968 14424 21974 14436
rect 22465 14433 22477 14436
rect 22511 14433 22523 14467
rect 22465 14427 22523 14433
rect 22741 14467 22799 14473
rect 22741 14433 22753 14467
rect 22787 14464 22799 14467
rect 22830 14464 22836 14476
rect 22787 14436 22836 14464
rect 22787 14433 22799 14436
rect 22741 14427 22799 14433
rect 22830 14424 22836 14436
rect 22888 14424 22894 14476
rect 24026 14424 24032 14476
rect 24084 14464 24090 14476
rect 25869 14467 25927 14473
rect 25869 14464 25881 14467
rect 24084 14436 25881 14464
rect 24084 14424 24090 14436
rect 25869 14433 25881 14436
rect 25915 14433 25927 14467
rect 25869 14427 25927 14433
rect 26145 14467 26203 14473
rect 26145 14433 26157 14467
rect 26191 14464 26203 14467
rect 26234 14464 26240 14476
rect 26191 14436 26240 14464
rect 26191 14433 26203 14436
rect 26145 14427 26203 14433
rect 26234 14424 26240 14436
rect 26292 14464 26298 14476
rect 27154 14464 27160 14476
rect 26292 14436 27160 14464
rect 26292 14424 26298 14436
rect 27154 14424 27160 14436
rect 27212 14424 27218 14476
rect 27522 14424 27528 14476
rect 27580 14464 27586 14476
rect 28169 14467 28227 14473
rect 28169 14464 28181 14467
rect 27580 14436 28181 14464
rect 27580 14424 27586 14436
rect 28169 14433 28181 14436
rect 28215 14433 28227 14467
rect 28169 14427 28227 14433
rect 19610 14356 19616 14408
rect 19668 14356 19674 14408
rect 22186 14356 22192 14408
rect 22244 14396 22250 14408
rect 25041 14399 25099 14405
rect 22244 14368 22324 14396
rect 22244 14356 22250 14368
rect 20901 14331 20959 14337
rect 20901 14297 20913 14331
rect 20947 14328 20959 14331
rect 21174 14328 21180 14340
rect 20947 14300 21180 14328
rect 20947 14297 20959 14300
rect 20901 14291 20959 14297
rect 21174 14288 21180 14300
rect 21232 14288 21238 14340
rect 22296 14328 22324 14368
rect 25041 14365 25053 14399
rect 25087 14396 25099 14399
rect 25222 14396 25228 14408
rect 25087 14368 25228 14396
rect 25087 14365 25099 14368
rect 25041 14359 25099 14365
rect 25222 14356 25228 14368
rect 25280 14356 25286 14408
rect 25314 14356 25320 14408
rect 25372 14396 25378 14408
rect 25685 14399 25743 14405
rect 25685 14396 25697 14399
rect 25372 14368 25697 14396
rect 25372 14356 25378 14368
rect 25685 14365 25697 14368
rect 25731 14365 25743 14399
rect 25685 14359 25743 14365
rect 22126 14300 22232 14328
rect 22296 14300 23230 14328
rect 19702 14220 19708 14272
rect 19760 14220 19766 14272
rect 22204 14260 22232 14300
rect 25406 14288 25412 14340
rect 25464 14288 25470 14340
rect 27338 14288 27344 14340
rect 27396 14288 27402 14340
rect 27890 14288 27896 14340
rect 27948 14288 27954 14340
rect 22278 14260 22284 14272
rect 22204 14232 22284 14260
rect 22278 14220 22284 14232
rect 22336 14260 22342 14272
rect 23658 14260 23664 14272
rect 22336 14232 23664 14260
rect 22336 14220 22342 14232
rect 23658 14220 23664 14232
rect 23716 14220 23722 14272
rect 24394 14220 24400 14272
rect 24452 14220 24458 14272
rect 25317 14263 25375 14269
rect 25317 14229 25329 14263
rect 25363 14260 25375 14263
rect 25424 14260 25452 14288
rect 25363 14232 25452 14260
rect 25363 14229 25375 14232
rect 25317 14223 25375 14229
rect 25774 14220 25780 14272
rect 25832 14220 25838 14272
rect 1104 14170 38824 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 35594 14170
rect 35646 14118 35658 14170
rect 35710 14118 35722 14170
rect 35774 14118 35786 14170
rect 35838 14118 35850 14170
rect 35902 14118 38824 14170
rect 1104 14096 38824 14118
rect 19702 14016 19708 14068
rect 19760 14056 19766 14068
rect 20441 14059 20499 14065
rect 20441 14056 20453 14059
rect 19760 14028 20453 14056
rect 19760 14016 19766 14028
rect 20441 14025 20453 14028
rect 20487 14025 20499 14059
rect 22278 14056 22284 14068
rect 20441 14019 20499 14025
rect 21652 14028 22284 14056
rect 18782 13948 18788 14000
rect 18840 13988 18846 14000
rect 18877 13991 18935 13997
rect 18877 13988 18889 13991
rect 18840 13960 18889 13988
rect 18840 13948 18846 13960
rect 18877 13957 18889 13960
rect 18923 13957 18935 13991
rect 20622 13988 20628 14000
rect 20102 13960 20628 13988
rect 18877 13951 18935 13957
rect 20622 13948 20628 13960
rect 20680 13988 20686 14000
rect 21652 13988 21680 14028
rect 22278 14016 22284 14028
rect 22336 14016 22342 14068
rect 25498 14056 25504 14068
rect 25148 14028 25504 14056
rect 20680 13960 21680 13988
rect 20680 13948 20686 13960
rect 21910 13948 21916 14000
rect 21968 13988 21974 14000
rect 21968 13960 22968 13988
rect 21968 13948 21974 13960
rect 20898 13880 20904 13932
rect 20956 13920 20962 13932
rect 22940 13929 22968 13960
rect 23658 13948 23664 14000
rect 23716 13948 23722 14000
rect 25148 13997 25176 14028
rect 25498 14016 25504 14028
rect 25556 14016 25562 14068
rect 25774 14016 25780 14068
rect 25832 14056 25838 14068
rect 26973 14059 27031 14065
rect 26973 14056 26985 14059
rect 25832 14028 26985 14056
rect 25832 14016 25838 14028
rect 26973 14025 26985 14028
rect 27019 14025 27031 14059
rect 26973 14019 27031 14025
rect 27890 14016 27896 14068
rect 27948 14016 27954 14068
rect 25133 13991 25191 13997
rect 25133 13957 25145 13991
rect 25179 13957 25191 13991
rect 26694 13988 26700 14000
rect 26358 13960 26700 13988
rect 25133 13951 25191 13957
rect 26694 13948 26700 13960
rect 26752 13948 26758 14000
rect 22005 13923 22063 13929
rect 22005 13920 22017 13923
rect 20956 13892 22017 13920
rect 20956 13880 20962 13892
rect 22005 13889 22017 13892
rect 22051 13889 22063 13923
rect 22005 13883 22063 13889
rect 22925 13923 22983 13929
rect 22925 13889 22937 13923
rect 22971 13889 22983 13923
rect 22925 13883 22983 13889
rect 27706 13880 27712 13932
rect 27764 13880 27770 13932
rect 18598 13812 18604 13864
rect 18656 13812 18662 13864
rect 20349 13855 20407 13861
rect 20349 13821 20361 13855
rect 20395 13852 20407 13855
rect 20993 13855 21051 13861
rect 20993 13852 21005 13855
rect 20395 13824 21005 13852
rect 20395 13821 20407 13824
rect 20349 13815 20407 13821
rect 20993 13821 21005 13824
rect 21039 13852 21051 13855
rect 21039 13824 21864 13852
rect 21039 13821 21051 13824
rect 20993 13815 21051 13821
rect 21836 13784 21864 13824
rect 21910 13812 21916 13864
rect 21968 13812 21974 13864
rect 23198 13812 23204 13864
rect 23256 13812 23262 13864
rect 24486 13812 24492 13864
rect 24544 13812 24550 13864
rect 24854 13812 24860 13864
rect 24912 13812 24918 13864
rect 25866 13812 25872 13864
rect 25924 13852 25930 13864
rect 26605 13855 26663 13861
rect 26605 13852 26617 13855
rect 25924 13824 26617 13852
rect 25924 13812 25930 13824
rect 26605 13821 26617 13824
rect 26651 13852 26663 13855
rect 27525 13855 27583 13861
rect 27525 13852 27537 13855
rect 26651 13824 27537 13852
rect 26651 13821 26663 13824
rect 26605 13815 26663 13821
rect 27525 13821 27537 13824
rect 27571 13821 27583 13855
rect 27525 13815 27583 13821
rect 21836 13756 22094 13784
rect 22066 13716 22094 13756
rect 22186 13716 22192 13728
rect 22066 13688 22192 13716
rect 22186 13676 22192 13688
rect 22244 13676 22250 13728
rect 22281 13719 22339 13725
rect 22281 13685 22293 13719
rect 22327 13716 22339 13719
rect 24504 13716 24532 13812
rect 22327 13688 24532 13716
rect 24673 13719 24731 13725
rect 22327 13685 22339 13688
rect 22281 13679 22339 13685
rect 24673 13685 24685 13719
rect 24719 13716 24731 13719
rect 25222 13716 25228 13728
rect 24719 13688 25228 13716
rect 24719 13685 24731 13688
rect 24673 13679 24731 13685
rect 25222 13676 25228 13688
rect 25280 13676 25286 13728
rect 1104 13626 38824 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38824 13626
rect 1104 13552 38824 13574
rect 10134 13472 10140 13524
rect 10192 13512 10198 13524
rect 19705 13515 19763 13521
rect 10192 13484 12434 13512
rect 10192 13472 10198 13484
rect 12406 13444 12434 13484
rect 19705 13481 19717 13515
rect 19751 13512 19763 13515
rect 21910 13512 21916 13524
rect 19751 13484 21916 13512
rect 19751 13481 19763 13484
rect 19705 13475 19763 13481
rect 21910 13472 21916 13484
rect 21968 13472 21974 13524
rect 23198 13472 23204 13524
rect 23256 13472 23262 13524
rect 24026 13472 24032 13524
rect 24084 13512 24090 13524
rect 27525 13515 27583 13521
rect 24084 13484 26234 13512
rect 24084 13472 24090 13484
rect 20809 13447 20867 13453
rect 12406 13416 20760 13444
rect 19521 13379 19579 13385
rect 19521 13345 19533 13379
rect 19567 13376 19579 13379
rect 19610 13376 19616 13388
rect 19567 13348 19616 13376
rect 19567 13345 19579 13348
rect 19521 13339 19579 13345
rect 19610 13336 19616 13348
rect 19668 13336 19674 13388
rect 20533 13379 20591 13385
rect 20533 13345 20545 13379
rect 20579 13345 20591 13379
rect 20732 13376 20760 13416
rect 20809 13413 20821 13447
rect 20855 13444 20867 13447
rect 20898 13444 20904 13456
rect 20855 13416 20904 13444
rect 20855 13413 20867 13416
rect 20809 13407 20867 13413
rect 20898 13404 20904 13416
rect 20956 13404 20962 13456
rect 23477 13447 23535 13453
rect 23477 13413 23489 13447
rect 23523 13413 23535 13447
rect 26206 13444 26234 13484
rect 27525 13481 27537 13515
rect 27571 13512 27583 13515
rect 27706 13512 27712 13524
rect 27571 13484 27712 13512
rect 27571 13481 27583 13484
rect 27525 13475 27583 13481
rect 27706 13472 27712 13484
rect 27764 13472 27770 13524
rect 23477 13407 23535 13413
rect 23952 13416 24256 13444
rect 26206 13416 28028 13444
rect 20732 13348 23060 13376
rect 20533 13339 20591 13345
rect 19426 13268 19432 13320
rect 19484 13268 19490 13320
rect 20441 13311 20499 13317
rect 20441 13308 20453 13311
rect 19996 13280 20453 13308
rect 19996 13184 20024 13280
rect 20441 13277 20453 13280
rect 20487 13277 20499 13311
rect 20441 13271 20499 13277
rect 19978 13132 19984 13184
rect 20036 13132 20042 13184
rect 20548 13172 20576 13339
rect 20714 13268 20720 13320
rect 20772 13308 20778 13320
rect 20901 13311 20959 13317
rect 20901 13308 20913 13311
rect 20772 13280 20913 13308
rect 20772 13268 20778 13280
rect 20901 13277 20913 13280
rect 20947 13277 20959 13311
rect 20901 13271 20959 13277
rect 22278 13268 22284 13320
rect 22336 13268 22342 13320
rect 21174 13200 21180 13252
rect 21232 13200 21238 13252
rect 22002 13172 22008 13184
rect 20548 13144 22008 13172
rect 22002 13132 22008 13144
rect 22060 13132 22066 13184
rect 22649 13175 22707 13181
rect 22649 13141 22661 13175
rect 22695 13172 22707 13175
rect 22922 13172 22928 13184
rect 22695 13144 22928 13172
rect 22695 13141 22707 13144
rect 22649 13135 22707 13141
rect 22922 13132 22928 13144
rect 22980 13132 22986 13184
rect 23032 13172 23060 13348
rect 23385 13311 23443 13317
rect 23385 13277 23397 13311
rect 23431 13308 23443 13311
rect 23492 13308 23520 13407
rect 23952 13376 23980 13416
rect 24228 13388 24256 13416
rect 23860 13348 23980 13376
rect 23860 13317 23888 13348
rect 24026 13336 24032 13388
rect 24084 13336 24090 13388
rect 24210 13336 24216 13388
rect 24268 13336 24274 13388
rect 24394 13336 24400 13388
rect 24452 13336 24458 13388
rect 24854 13336 24860 13388
rect 24912 13376 24918 13388
rect 28000 13385 28028 13416
rect 26973 13379 27031 13385
rect 24912 13348 26740 13376
rect 24912 13336 24918 13348
rect 23431 13280 23520 13308
rect 23845 13311 23903 13317
rect 23431 13277 23443 13280
rect 23385 13271 23443 13277
rect 23845 13277 23857 13311
rect 23891 13277 23903 13311
rect 23845 13271 23903 13277
rect 23937 13311 23995 13317
rect 23937 13277 23949 13311
rect 23983 13308 23995 13311
rect 24412 13308 24440 13336
rect 23983 13280 24440 13308
rect 25225 13311 25283 13317
rect 23983 13277 23995 13280
rect 23937 13271 23995 13277
rect 25225 13277 25237 13311
rect 25271 13308 25283 13311
rect 25314 13308 25320 13320
rect 25271 13280 25320 13308
rect 25271 13277 25283 13280
rect 25225 13271 25283 13277
rect 25314 13268 25320 13280
rect 25372 13268 25378 13320
rect 26712 13308 26740 13348
rect 26973 13345 26985 13379
rect 27019 13376 27031 13379
rect 27985 13379 28043 13385
rect 27019 13348 27844 13376
rect 27019 13345 27031 13348
rect 26973 13339 27031 13345
rect 27522 13308 27528 13320
rect 26712 13280 27528 13308
rect 27522 13268 27528 13280
rect 27580 13268 27586 13320
rect 27709 13311 27767 13317
rect 27709 13277 27721 13311
rect 27755 13277 27767 13311
rect 27816 13308 27844 13348
rect 27985 13345 27997 13379
rect 28031 13345 28043 13379
rect 27985 13339 28043 13345
rect 28074 13308 28080 13320
rect 27816 13280 28080 13308
rect 27709 13271 27767 13277
rect 26234 13200 26240 13252
rect 26292 13200 26298 13252
rect 27154 13200 27160 13252
rect 27212 13200 27218 13252
rect 26602 13172 26608 13184
rect 23032 13144 26608 13172
rect 26602 13132 26608 13144
rect 26660 13181 26666 13184
rect 26660 13175 26709 13181
rect 26660 13141 26663 13175
rect 26697 13141 26709 13175
rect 26660 13135 26709 13141
rect 27065 13175 27123 13181
rect 27065 13141 27077 13175
rect 27111 13172 27123 13175
rect 27724 13172 27752 13271
rect 28074 13268 28080 13280
rect 28132 13268 28138 13320
rect 29914 13172 29920 13184
rect 27111 13144 29920 13172
rect 27111 13141 27123 13144
rect 27065 13135 27123 13141
rect 26660 13132 26666 13135
rect 29914 13132 29920 13144
rect 29972 13132 29978 13184
rect 1104 13082 38824 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 35594 13082
rect 35646 13030 35658 13082
rect 35710 13030 35722 13082
rect 35774 13030 35786 13082
rect 35838 13030 35850 13082
rect 35902 13030 38824 13082
rect 1104 13008 38824 13030
rect 21174 12928 21180 12980
rect 21232 12968 21238 12980
rect 21269 12971 21327 12977
rect 21269 12968 21281 12971
rect 21232 12940 21281 12968
rect 21232 12928 21238 12940
rect 21269 12937 21281 12940
rect 21315 12937 21327 12971
rect 21269 12931 21327 12937
rect 22186 12928 22192 12980
rect 22244 12968 22250 12980
rect 22244 12940 23612 12968
rect 22244 12928 22250 12940
rect 19797 12903 19855 12909
rect 19797 12900 19809 12903
rect 6886 12872 19809 12900
rect 1394 12792 1400 12844
rect 1452 12792 1458 12844
rect 1581 12631 1639 12637
rect 1581 12597 1593 12631
rect 1627 12628 1639 12631
rect 6886 12628 6914 12872
rect 19797 12869 19809 12872
rect 19843 12900 19855 12903
rect 19978 12900 19984 12912
rect 19843 12872 19984 12900
rect 19843 12869 19855 12872
rect 19797 12863 19855 12869
rect 19978 12860 19984 12872
rect 20036 12860 20042 12912
rect 19153 12835 19211 12841
rect 19153 12801 19165 12835
rect 19199 12832 19211 12835
rect 19889 12835 19947 12841
rect 19199 12804 19472 12832
rect 19199 12801 19211 12804
rect 19153 12795 19211 12801
rect 19444 12705 19472 12804
rect 19889 12801 19901 12835
rect 19935 12832 19947 12835
rect 20441 12835 20499 12841
rect 20441 12832 20453 12835
rect 19935 12804 20453 12832
rect 19935 12801 19947 12804
rect 19889 12795 19947 12801
rect 20441 12801 20453 12804
rect 20487 12801 20499 12835
rect 20441 12795 20499 12801
rect 21450 12792 21456 12844
rect 21508 12792 21514 12844
rect 22830 12792 22836 12844
rect 22888 12841 22894 12844
rect 22888 12835 22916 12841
rect 22904 12801 22916 12835
rect 22888 12795 22916 12801
rect 22888 12792 22894 12795
rect 20070 12724 20076 12776
rect 20128 12724 20134 12776
rect 21082 12724 21088 12776
rect 21140 12764 21146 12776
rect 21821 12767 21879 12773
rect 21821 12764 21833 12767
rect 21140 12736 21833 12764
rect 21140 12724 21146 12736
rect 21821 12733 21833 12736
rect 21867 12733 21879 12767
rect 21821 12727 21879 12733
rect 22005 12767 22063 12773
rect 22005 12733 22017 12767
rect 22051 12733 22063 12767
rect 22005 12727 22063 12733
rect 19429 12699 19487 12705
rect 19429 12665 19441 12699
rect 19475 12665 19487 12699
rect 19429 12659 19487 12665
rect 1627 12600 6914 12628
rect 19337 12631 19395 12637
rect 1627 12597 1639 12600
rect 1581 12591 1639 12597
rect 19337 12597 19349 12631
rect 19383 12628 19395 12631
rect 19518 12628 19524 12640
rect 19383 12600 19524 12628
rect 19383 12597 19395 12600
rect 19337 12591 19395 12597
rect 19518 12588 19524 12600
rect 19576 12588 19582 12640
rect 22020 12628 22048 12727
rect 22370 12724 22376 12776
rect 22428 12764 22434 12776
rect 22741 12767 22799 12773
rect 22741 12764 22753 12767
rect 22428 12736 22753 12764
rect 22428 12724 22434 12736
rect 22741 12733 22753 12736
rect 22787 12733 22799 12767
rect 22741 12727 22799 12733
rect 23017 12767 23075 12773
rect 23017 12733 23029 12767
rect 23063 12764 23075 12767
rect 23198 12764 23204 12776
rect 23063 12736 23204 12764
rect 23063 12733 23075 12736
rect 23017 12727 23075 12733
rect 23198 12724 23204 12736
rect 23256 12764 23262 12776
rect 23584 12764 23612 12940
rect 26234 12928 26240 12980
rect 26292 12968 26298 12980
rect 27338 12968 27344 12980
rect 26292 12940 27344 12968
rect 26292 12928 26298 12940
rect 27338 12928 27344 12940
rect 27396 12968 27402 12980
rect 27396 12940 28856 12968
rect 27396 12928 27402 12940
rect 25884 12872 26372 12900
rect 24394 12792 24400 12844
rect 24452 12792 24458 12844
rect 25222 12792 25228 12844
rect 25280 12832 25286 12844
rect 25884 12841 25912 12872
rect 25409 12835 25467 12841
rect 25409 12832 25421 12835
rect 25280 12804 25421 12832
rect 25280 12792 25286 12804
rect 25409 12801 25421 12804
rect 25455 12801 25467 12835
rect 25409 12795 25467 12801
rect 25685 12835 25743 12841
rect 25685 12801 25697 12835
rect 25731 12801 25743 12835
rect 25685 12795 25743 12801
rect 25869 12835 25927 12841
rect 25869 12801 25881 12835
rect 25915 12801 25927 12835
rect 25869 12795 25927 12801
rect 26053 12835 26111 12841
rect 26053 12801 26065 12835
rect 26099 12801 26111 12835
rect 26053 12795 26111 12801
rect 24535 12767 24593 12773
rect 24535 12764 24547 12767
rect 23256 12736 23520 12764
rect 23584 12736 24547 12764
rect 23256 12724 23262 12736
rect 22465 12699 22523 12705
rect 22465 12665 22477 12699
rect 22511 12696 22523 12699
rect 22554 12696 22560 12708
rect 22511 12668 22560 12696
rect 22511 12665 22523 12668
rect 22465 12659 22523 12665
rect 22554 12656 22560 12668
rect 22612 12656 22618 12708
rect 23492 12696 23520 12736
rect 24535 12733 24547 12736
rect 24581 12733 24593 12767
rect 24535 12727 24593 12733
rect 24670 12724 24676 12776
rect 24728 12724 24734 12776
rect 25038 12724 25044 12776
rect 25096 12764 25102 12776
rect 25593 12767 25651 12773
rect 25593 12764 25605 12767
rect 25096 12736 25605 12764
rect 25096 12724 25102 12736
rect 25593 12733 25605 12736
rect 25639 12733 25651 12767
rect 25700 12764 25728 12795
rect 25958 12764 25964 12776
rect 25700 12736 25964 12764
rect 25593 12727 25651 12733
rect 25958 12724 25964 12736
rect 26016 12724 26022 12776
rect 23492 12668 24072 12696
rect 22922 12628 22928 12640
rect 22020 12600 22928 12628
rect 22922 12588 22928 12600
rect 22980 12588 22986 12640
rect 23658 12588 23664 12640
rect 23716 12588 23722 12640
rect 23750 12588 23756 12640
rect 23808 12588 23814 12640
rect 24044 12628 24072 12668
rect 24946 12656 24952 12708
rect 25004 12656 25010 12708
rect 25498 12656 25504 12708
rect 25556 12696 25562 12708
rect 26068 12696 26096 12795
rect 26234 12724 26240 12776
rect 26292 12724 26298 12776
rect 26344 12708 26372 12872
rect 28828 12844 28856 12940
rect 26605 12835 26663 12841
rect 26605 12832 26617 12835
rect 26436 12804 26617 12832
rect 26436 12776 26464 12804
rect 26605 12801 26617 12804
rect 26651 12801 26663 12835
rect 26605 12795 26663 12801
rect 26786 12792 26792 12844
rect 26844 12792 26850 12844
rect 28810 12792 28816 12844
rect 28868 12792 28874 12844
rect 26418 12724 26424 12776
rect 26476 12724 26482 12776
rect 27433 12767 27491 12773
rect 27433 12733 27445 12767
rect 27479 12764 27491 12767
rect 27479 12736 27568 12764
rect 27479 12733 27491 12736
rect 27433 12727 27491 12733
rect 25556 12668 26096 12696
rect 25556 12656 25562 12668
rect 26326 12656 26332 12708
rect 26384 12696 26390 12708
rect 26513 12699 26571 12705
rect 26513 12696 26525 12699
rect 26384 12668 26525 12696
rect 26384 12656 26390 12668
rect 26513 12665 26525 12668
rect 26559 12665 26571 12699
rect 26513 12659 26571 12665
rect 27540 12640 27568 12736
rect 27706 12724 27712 12776
rect 27764 12724 27770 12776
rect 29457 12767 29515 12773
rect 29457 12733 29469 12767
rect 29503 12764 29515 12767
rect 29546 12764 29552 12776
rect 29503 12736 29552 12764
rect 29503 12733 29515 12736
rect 29457 12727 29515 12733
rect 29546 12724 29552 12736
rect 29604 12724 29610 12776
rect 24394 12628 24400 12640
rect 24044 12600 24400 12628
rect 24394 12588 24400 12600
rect 24452 12588 24458 12640
rect 24486 12588 24492 12640
rect 24544 12628 24550 12640
rect 25777 12631 25835 12637
rect 25777 12628 25789 12631
rect 24544 12600 25789 12628
rect 24544 12588 24550 12600
rect 25777 12597 25789 12600
rect 25823 12597 25835 12631
rect 25777 12591 25835 12597
rect 27522 12588 27528 12640
rect 27580 12588 27586 12640
rect 1104 12538 38824 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38824 12538
rect 1104 12464 38824 12486
rect 19978 12424 19984 12436
rect 18984 12396 19984 12424
rect 18598 12248 18604 12300
rect 18656 12248 18662 12300
rect 18984 12297 19012 12396
rect 19978 12384 19984 12396
rect 20036 12424 20042 12436
rect 20993 12427 21051 12433
rect 20036 12396 20944 12424
rect 20036 12384 20042 12396
rect 18969 12291 19027 12297
rect 18969 12257 18981 12291
rect 19015 12257 19027 12291
rect 20806 12288 20812 12300
rect 18969 12251 19027 12257
rect 19260 12260 20812 12288
rect 18049 12223 18107 12229
rect 18049 12189 18061 12223
rect 18095 12220 18107 12223
rect 18616 12220 18644 12248
rect 19260 12229 19288 12260
rect 20806 12248 20812 12260
rect 20864 12248 20870 12300
rect 20916 12288 20944 12396
rect 20993 12393 21005 12427
rect 21039 12424 21051 12427
rect 21082 12424 21088 12436
rect 21039 12396 21088 12424
rect 21039 12393 21051 12396
rect 20993 12387 21051 12393
rect 21082 12384 21088 12396
rect 21140 12384 21146 12436
rect 21450 12384 21456 12436
rect 21508 12424 21514 12436
rect 21545 12427 21603 12433
rect 21545 12424 21557 12427
rect 21508 12396 21557 12424
rect 21508 12384 21514 12396
rect 21545 12393 21557 12396
rect 21591 12393 21603 12427
rect 21545 12387 21603 12393
rect 23658 12384 23664 12436
rect 23716 12424 23722 12436
rect 24581 12427 24639 12433
rect 24581 12424 24593 12427
rect 23716 12396 24593 12424
rect 23716 12384 23722 12396
rect 24581 12393 24593 12396
rect 24627 12393 24639 12427
rect 24581 12387 24639 12393
rect 27706 12384 27712 12436
rect 27764 12424 27770 12436
rect 27985 12427 28043 12433
rect 27985 12424 27997 12427
rect 27764 12396 27997 12424
rect 27764 12384 27770 12396
rect 27985 12393 27997 12396
rect 28031 12393 28043 12427
rect 27985 12387 28043 12393
rect 26418 12356 26424 12368
rect 26160 12328 26424 12356
rect 22097 12291 22155 12297
rect 22097 12288 22109 12291
rect 20916 12260 22109 12288
rect 22097 12257 22109 12260
rect 22143 12257 22155 12291
rect 22097 12251 22155 12257
rect 22922 12248 22928 12300
rect 22980 12248 22986 12300
rect 24213 12291 24271 12297
rect 24213 12257 24225 12291
rect 24259 12288 24271 12291
rect 24259 12260 25636 12288
rect 24259 12257 24271 12260
rect 24213 12251 24271 12257
rect 19245 12223 19303 12229
rect 19245 12220 19257 12223
rect 18095 12192 18368 12220
rect 18616 12192 19257 12220
rect 18095 12189 18107 12192
rect 18049 12183 18107 12189
rect 18230 12044 18236 12096
rect 18288 12044 18294 12096
rect 18340 12093 18368 12192
rect 19245 12189 19257 12192
rect 19291 12189 19303 12223
rect 19245 12183 19303 12189
rect 20622 12180 20628 12232
rect 20680 12180 20686 12232
rect 21913 12223 21971 12229
rect 21913 12189 21925 12223
rect 21959 12220 21971 12223
rect 22002 12220 22008 12232
rect 21959 12192 22008 12220
rect 21959 12189 21971 12192
rect 21913 12183 21971 12189
rect 22002 12180 22008 12192
rect 22060 12180 22066 12232
rect 23842 12180 23848 12232
rect 23900 12180 23906 12232
rect 24029 12223 24087 12229
rect 24029 12189 24041 12223
rect 24075 12220 24087 12223
rect 24489 12223 24547 12229
rect 24489 12220 24501 12223
rect 24075 12192 24501 12220
rect 24075 12189 24087 12192
rect 24029 12183 24087 12189
rect 24489 12189 24501 12192
rect 24535 12220 24547 12223
rect 24535 12192 24624 12220
rect 24535 12189 24547 12192
rect 24489 12183 24547 12189
rect 19426 12152 19432 12164
rect 18708 12124 19432 12152
rect 18708 12096 18736 12124
rect 19426 12112 19432 12124
rect 19484 12112 19490 12164
rect 19518 12112 19524 12164
rect 19576 12112 19582 12164
rect 24596 12096 24624 12192
rect 25406 12180 25412 12232
rect 25464 12180 25470 12232
rect 25608 12229 25636 12260
rect 25866 12248 25872 12300
rect 25924 12248 25930 12300
rect 26160 12297 26188 12328
rect 26418 12316 26424 12328
rect 26476 12356 26482 12368
rect 29546 12356 29552 12368
rect 26476 12328 29552 12356
rect 26476 12316 26482 12328
rect 26145 12291 26203 12297
rect 26145 12257 26157 12291
rect 26191 12257 26203 12291
rect 26145 12251 26203 12257
rect 26602 12248 26608 12300
rect 26660 12248 26666 12300
rect 27264 12288 27292 12328
rect 29546 12316 29552 12328
rect 29604 12316 29610 12368
rect 27080 12260 27292 12288
rect 27433 12291 27491 12297
rect 25593 12223 25651 12229
rect 25593 12189 25605 12223
rect 25639 12189 25651 12223
rect 25593 12183 25651 12189
rect 25958 12180 25964 12232
rect 26016 12220 26022 12232
rect 26234 12220 26240 12232
rect 26016 12192 26240 12220
rect 26016 12180 26022 12192
rect 26234 12180 26240 12192
rect 26292 12180 26298 12232
rect 26878 12180 26884 12232
rect 26936 12180 26942 12232
rect 26970 12180 26976 12232
rect 27028 12220 27034 12232
rect 27080 12229 27108 12260
rect 27433 12257 27445 12291
rect 27479 12288 27491 12291
rect 28074 12288 28080 12300
rect 27479 12260 28080 12288
rect 27479 12257 27491 12260
rect 27433 12251 27491 12257
rect 28074 12248 28080 12260
rect 28132 12288 28138 12300
rect 28132 12260 28764 12288
rect 28132 12248 28138 12260
rect 28736 12232 28764 12260
rect 27065 12223 27123 12229
rect 27065 12220 27077 12223
rect 27028 12192 27077 12220
rect 27028 12180 27034 12192
rect 27065 12189 27077 12192
rect 27111 12189 27123 12223
rect 27065 12183 27123 12189
rect 27246 12180 27252 12232
rect 27304 12180 27310 12232
rect 27709 12223 27767 12229
rect 27709 12189 27721 12223
rect 27755 12189 27767 12223
rect 27709 12183 27767 12189
rect 25501 12155 25559 12161
rect 25501 12152 25513 12155
rect 24964 12124 25513 12152
rect 18325 12087 18383 12093
rect 18325 12053 18337 12087
rect 18371 12053 18383 12087
rect 18325 12047 18383 12053
rect 18690 12044 18696 12096
rect 18748 12044 18754 12096
rect 18782 12044 18788 12096
rect 18840 12044 18846 12096
rect 22005 12087 22063 12093
rect 22005 12053 22017 12087
rect 22051 12084 22063 12087
rect 22373 12087 22431 12093
rect 22373 12084 22385 12087
rect 22051 12056 22385 12084
rect 22051 12053 22063 12056
rect 22005 12047 22063 12053
rect 22373 12053 22385 12056
rect 22419 12053 22431 12087
rect 22373 12047 22431 12053
rect 24578 12044 24584 12096
rect 24636 12044 24642 12096
rect 24964 12093 24992 12124
rect 25501 12121 25513 12124
rect 25547 12121 25559 12155
rect 25501 12115 25559 12121
rect 25731 12155 25789 12161
rect 25731 12121 25743 12155
rect 25777 12152 25789 12155
rect 26418 12152 26424 12164
rect 25777 12124 26424 12152
rect 25777 12121 25789 12124
rect 25731 12115 25789 12121
rect 26418 12112 26424 12124
rect 26476 12112 26482 12164
rect 26513 12155 26571 12161
rect 26513 12121 26525 12155
rect 26559 12152 26571 12155
rect 26896 12152 26924 12180
rect 27724 12152 27752 12183
rect 28166 12180 28172 12232
rect 28224 12180 28230 12232
rect 28718 12180 28724 12232
rect 28776 12180 28782 12232
rect 26559 12124 29776 12152
rect 26559 12121 26571 12124
rect 26513 12115 26571 12121
rect 29748 12096 29776 12124
rect 24949 12087 25007 12093
rect 24949 12053 24961 12087
rect 24995 12053 25007 12087
rect 24949 12047 25007 12053
rect 25222 12044 25228 12096
rect 25280 12044 25286 12096
rect 25958 12044 25964 12096
rect 26016 12044 26022 12096
rect 27614 12044 27620 12096
rect 27672 12044 27678 12096
rect 29730 12044 29736 12096
rect 29788 12044 29794 12096
rect 1104 11994 38824 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 35594 11994
rect 35646 11942 35658 11994
rect 35710 11942 35722 11994
rect 35774 11942 35786 11994
rect 35838 11942 35850 11994
rect 35902 11942 38824 11994
rect 1104 11920 38824 11942
rect 18230 11840 18236 11892
rect 18288 11840 18294 11892
rect 18598 11840 18604 11892
rect 18656 11840 18662 11892
rect 20438 11840 20444 11892
rect 20496 11840 20502 11892
rect 22281 11883 22339 11889
rect 22281 11849 22293 11883
rect 22327 11880 22339 11883
rect 22327 11852 24716 11880
rect 22327 11849 22339 11852
rect 22281 11843 22339 11849
rect 18248 11676 18276 11840
rect 18616 11744 18644 11840
rect 24688 11824 24716 11852
rect 26418 11840 26424 11892
rect 26476 11840 26482 11892
rect 26789 11883 26847 11889
rect 26789 11849 26801 11883
rect 26835 11880 26847 11883
rect 28166 11880 28172 11892
rect 26835 11852 28172 11880
rect 26835 11849 26847 11852
rect 26789 11843 26847 11849
rect 28166 11840 28172 11852
rect 28224 11840 28230 11892
rect 20533 11815 20591 11821
rect 20533 11812 20545 11815
rect 20194 11784 20545 11812
rect 20533 11781 20545 11784
rect 20579 11812 20591 11815
rect 20622 11812 20628 11824
rect 20579 11784 20628 11812
rect 20579 11781 20591 11784
rect 20533 11775 20591 11781
rect 20622 11772 20628 11784
rect 20680 11772 20686 11824
rect 20901 11815 20959 11821
rect 20901 11781 20913 11815
rect 20947 11812 20959 11815
rect 22094 11812 22100 11824
rect 20947 11784 22100 11812
rect 20947 11781 20959 11784
rect 20901 11775 20959 11781
rect 22094 11772 22100 11784
rect 22152 11772 22158 11824
rect 23198 11812 23204 11824
rect 22848 11784 23204 11812
rect 18693 11747 18751 11753
rect 18693 11744 18705 11747
rect 18616 11716 18705 11744
rect 18693 11713 18705 11716
rect 18739 11713 18751 11747
rect 18693 11707 18751 11713
rect 22186 11704 22192 11756
rect 22244 11704 22250 11756
rect 22848 11753 22876 11784
rect 23198 11772 23204 11784
rect 23256 11772 23262 11824
rect 23566 11772 23572 11824
rect 23624 11812 23630 11824
rect 23624 11784 23782 11812
rect 23624 11772 23630 11784
rect 24670 11772 24676 11824
rect 24728 11812 24734 11824
rect 25869 11815 25927 11821
rect 25869 11812 25881 11815
rect 24728 11784 25881 11812
rect 24728 11772 24734 11784
rect 25869 11781 25881 11784
rect 25915 11781 25927 11815
rect 26436 11812 26464 11840
rect 26973 11815 27031 11821
rect 26973 11812 26985 11815
rect 26436 11784 26985 11812
rect 25869 11775 25927 11781
rect 26973 11781 26985 11784
rect 27019 11781 27031 11815
rect 26973 11775 27031 11781
rect 22649 11747 22707 11753
rect 22649 11713 22661 11747
rect 22695 11744 22707 11747
rect 22833 11747 22891 11753
rect 22695 11716 22784 11744
rect 22695 11713 22707 11716
rect 22649 11707 22707 11713
rect 18969 11679 19027 11685
rect 18969 11676 18981 11679
rect 18248 11648 18981 11676
rect 18969 11645 18981 11648
rect 19015 11645 19027 11679
rect 18969 11639 19027 11645
rect 22465 11679 22523 11685
rect 22465 11645 22477 11679
rect 22511 11676 22523 11679
rect 22554 11676 22560 11688
rect 22511 11648 22560 11676
rect 22511 11645 22523 11648
rect 22465 11639 22523 11645
rect 22554 11636 22560 11648
rect 22612 11676 22618 11688
rect 22756 11676 22784 11716
rect 22833 11713 22845 11747
rect 22879 11713 22891 11747
rect 22833 11707 22891 11713
rect 25130 11704 25136 11756
rect 25188 11744 25194 11756
rect 25593 11747 25651 11753
rect 25593 11744 25605 11747
rect 25188 11716 25605 11744
rect 25188 11704 25194 11716
rect 25593 11713 25605 11716
rect 25639 11713 25651 11747
rect 26326 11744 26332 11756
rect 25593 11707 25651 11713
rect 25884 11716 26332 11744
rect 22922 11676 22928 11688
rect 22612 11648 22928 11676
rect 22612 11636 22618 11648
rect 22922 11636 22928 11648
rect 22980 11636 22986 11688
rect 23017 11679 23075 11685
rect 23017 11645 23029 11679
rect 23063 11645 23075 11679
rect 23017 11639 23075 11645
rect 23293 11679 23351 11685
rect 23293 11645 23305 11679
rect 23339 11676 23351 11679
rect 23750 11676 23756 11688
rect 23339 11648 23756 11676
rect 23339 11645 23351 11648
rect 23293 11639 23351 11645
rect 20806 11568 20812 11620
rect 20864 11608 20870 11620
rect 23032 11608 23060 11639
rect 23750 11636 23756 11648
rect 23808 11636 23814 11688
rect 25884 11685 25912 11716
rect 26326 11704 26332 11716
rect 26384 11704 26390 11756
rect 26421 11747 26479 11753
rect 26421 11713 26433 11747
rect 26467 11744 26479 11747
rect 26878 11744 26884 11756
rect 26467 11716 26884 11744
rect 26467 11713 26479 11716
rect 26421 11707 26479 11713
rect 26878 11704 26884 11716
rect 26936 11744 26942 11756
rect 27137 11745 27195 11751
rect 26936 11742 27016 11744
rect 27137 11742 27149 11745
rect 26936 11716 27149 11742
rect 26936 11704 26942 11716
rect 26988 11714 27149 11716
rect 27137 11711 27149 11714
rect 27183 11711 27195 11745
rect 27137 11705 27195 11711
rect 28810 11704 28816 11756
rect 28868 11744 28874 11756
rect 28868 11716 28934 11744
rect 28868 11704 28874 11716
rect 29638 11704 29644 11756
rect 29696 11704 29702 11756
rect 25409 11679 25467 11685
rect 25409 11676 25421 11679
rect 24780 11648 25421 11676
rect 20864 11580 23060 11608
rect 20864 11568 20870 11580
rect 21818 11500 21824 11552
rect 21876 11500 21882 11552
rect 22741 11543 22799 11549
rect 22741 11509 22753 11543
rect 22787 11540 22799 11543
rect 23106 11540 23112 11552
rect 22787 11512 23112 11540
rect 22787 11509 22799 11512
rect 22741 11503 22799 11509
rect 23106 11500 23112 11512
rect 23164 11500 23170 11552
rect 24578 11500 24584 11552
rect 24636 11540 24642 11552
rect 24780 11549 24808 11648
rect 25409 11645 25421 11648
rect 25455 11645 25467 11679
rect 25869 11679 25927 11685
rect 25869 11676 25881 11679
rect 25409 11639 25467 11645
rect 25608 11648 25881 11676
rect 25608 11620 25636 11648
rect 25869 11645 25881 11648
rect 25915 11645 25927 11679
rect 25869 11639 25927 11645
rect 26237 11679 26295 11685
rect 26237 11645 26249 11679
rect 26283 11676 26295 11679
rect 27341 11679 27399 11685
rect 27341 11676 27353 11679
rect 26283 11648 26464 11676
rect 26283 11645 26295 11648
rect 26237 11639 26295 11645
rect 25590 11568 25596 11620
rect 25648 11568 25654 11620
rect 26436 11552 26464 11648
rect 26620 11648 27353 11676
rect 26620 11552 26648 11648
rect 27341 11645 27353 11648
rect 27387 11645 27399 11679
rect 27341 11639 27399 11645
rect 27356 11608 27384 11639
rect 27522 11636 27528 11688
rect 27580 11636 27586 11688
rect 27798 11636 27804 11688
rect 27856 11636 27862 11688
rect 29549 11679 29607 11685
rect 29549 11645 29561 11679
rect 29595 11676 29607 11679
rect 29595 11648 29776 11676
rect 29595 11645 29607 11648
rect 29549 11639 29607 11645
rect 27356 11580 27660 11608
rect 27632 11552 27660 11580
rect 29748 11552 29776 11648
rect 29914 11568 29920 11620
rect 29972 11608 29978 11620
rect 38194 11608 38200 11620
rect 29972 11580 38200 11608
rect 29972 11568 29978 11580
rect 38194 11568 38200 11580
rect 38252 11568 38258 11620
rect 24765 11543 24823 11549
rect 24765 11540 24777 11543
rect 24636 11512 24777 11540
rect 24636 11500 24642 11512
rect 24765 11509 24777 11512
rect 24811 11509 24823 11543
rect 24765 11503 24823 11509
rect 24854 11500 24860 11552
rect 24912 11500 24918 11552
rect 25038 11500 25044 11552
rect 25096 11540 25102 11552
rect 25685 11543 25743 11549
rect 25685 11540 25697 11543
rect 25096 11512 25697 11540
rect 25096 11500 25102 11512
rect 25685 11509 25697 11512
rect 25731 11509 25743 11543
rect 25685 11503 25743 11509
rect 26418 11500 26424 11552
rect 26476 11500 26482 11552
rect 26602 11500 26608 11552
rect 26660 11500 26666 11552
rect 27614 11500 27620 11552
rect 27672 11500 27678 11552
rect 29730 11500 29736 11552
rect 29788 11500 29794 11552
rect 29822 11500 29828 11552
rect 29880 11500 29886 11552
rect 1104 11450 38824 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38824 11450
rect 1104 11376 38824 11398
rect 18782 11296 18788 11348
rect 18840 11336 18846 11348
rect 19613 11339 19671 11345
rect 19613 11336 19625 11339
rect 18840 11308 19625 11336
rect 18840 11296 18846 11308
rect 19613 11305 19625 11308
rect 19659 11305 19671 11339
rect 19613 11299 19671 11305
rect 20806 11296 20812 11348
rect 20864 11296 20870 11348
rect 22094 11296 22100 11348
rect 22152 11336 22158 11348
rect 23014 11336 23020 11348
rect 22152 11308 23020 11336
rect 22152 11296 22158 11308
rect 23014 11296 23020 11308
rect 23072 11296 23078 11348
rect 25222 11296 25228 11348
rect 25280 11296 25286 11348
rect 25314 11296 25320 11348
rect 25372 11336 25378 11348
rect 25409 11339 25467 11345
rect 25409 11336 25421 11339
rect 25372 11308 25421 11336
rect 25372 11296 25378 11308
rect 25409 11305 25421 11308
rect 25455 11305 25467 11339
rect 25409 11299 25467 11305
rect 25958 11296 25964 11348
rect 26016 11296 26022 11348
rect 26142 11296 26148 11348
rect 26200 11336 26206 11348
rect 26237 11339 26295 11345
rect 26237 11336 26249 11339
rect 26200 11308 26249 11336
rect 26200 11296 26206 11308
rect 26237 11305 26249 11308
rect 26283 11336 26295 11339
rect 26878 11336 26884 11348
rect 26283 11308 26884 11336
rect 26283 11305 26295 11308
rect 26237 11299 26295 11305
rect 26878 11296 26884 11308
rect 26936 11296 26942 11348
rect 27798 11296 27804 11348
rect 27856 11296 27862 11348
rect 27890 11296 27896 11348
rect 27948 11296 27954 11348
rect 29089 11339 29147 11345
rect 29089 11305 29101 11339
rect 29135 11336 29147 11339
rect 29546 11336 29552 11348
rect 29135 11308 29552 11336
rect 29135 11305 29147 11308
rect 29089 11299 29147 11305
rect 29546 11296 29552 11308
rect 29604 11296 29610 11348
rect 29822 11296 29828 11348
rect 29880 11296 29886 11348
rect 20257 11203 20315 11209
rect 20257 11169 20269 11203
rect 20303 11200 20315 11203
rect 20438 11200 20444 11212
rect 20303 11172 20444 11200
rect 20303 11169 20315 11172
rect 20257 11163 20315 11169
rect 20438 11160 20444 11172
rect 20496 11160 20502 11212
rect 20717 11203 20775 11209
rect 20717 11169 20729 11203
rect 20763 11200 20775 11203
rect 20824 11200 20852 11296
rect 23198 11228 23204 11280
rect 23256 11268 23262 11280
rect 23566 11268 23572 11280
rect 23256 11240 23572 11268
rect 23256 11228 23262 11240
rect 23566 11228 23572 11240
rect 23624 11268 23630 11280
rect 23624 11240 24164 11268
rect 23624 11228 23630 11240
rect 20763 11172 20852 11200
rect 20763 11169 20775 11172
rect 20717 11163 20775 11169
rect 22186 11160 22192 11212
rect 22244 11200 22250 11212
rect 24136 11209 24164 11240
rect 24121 11203 24179 11209
rect 22244 11172 23888 11200
rect 22244 11160 22250 11172
rect 20622 11092 20628 11144
rect 20680 11092 20686 11144
rect 23124 11141 23152 11172
rect 23860 11144 23888 11172
rect 24121 11169 24133 11203
rect 24167 11169 24179 11203
rect 24121 11163 24179 11169
rect 23017 11135 23075 11141
rect 23017 11101 23029 11135
rect 23063 11101 23075 11135
rect 23017 11095 23075 11101
rect 23109 11135 23167 11141
rect 23109 11101 23121 11135
rect 23155 11101 23167 11135
rect 23109 11095 23167 11101
rect 23477 11135 23535 11141
rect 23477 11101 23489 11135
rect 23523 11132 23535 11135
rect 23569 11135 23627 11141
rect 23569 11132 23581 11135
rect 23523 11104 23581 11132
rect 23523 11101 23535 11104
rect 23477 11095 23535 11101
rect 23569 11101 23581 11104
rect 23615 11101 23627 11135
rect 23569 11095 23627 11101
rect 20640 10996 20668 11092
rect 20990 11024 20996 11076
rect 21048 11024 21054 11076
rect 22741 11067 22799 11073
rect 21376 11036 21482 11064
rect 21376 10996 21404 11036
rect 22741 11033 22753 11067
rect 22787 11064 22799 11067
rect 22922 11064 22928 11076
rect 22787 11036 22928 11064
rect 22787 11033 22799 11036
rect 22741 11027 22799 11033
rect 22922 11024 22928 11036
rect 22980 11024 22986 11076
rect 20640 10968 21404 10996
rect 22830 10956 22836 11008
rect 22888 10956 22894 11008
rect 23032 10996 23060 11095
rect 23842 11092 23848 11144
rect 23900 11092 23906 11144
rect 24136 11132 24164 11163
rect 25130 11160 25136 11212
rect 25188 11160 25194 11212
rect 25240 11200 25268 11296
rect 25593 11203 25651 11209
rect 25593 11200 25605 11203
rect 25240 11172 25605 11200
rect 25593 11169 25605 11172
rect 25639 11169 25651 11203
rect 25593 11163 25651 11169
rect 25869 11203 25927 11209
rect 25869 11169 25881 11203
rect 25915 11200 25927 11203
rect 25976 11200 26004 11296
rect 26602 11268 26608 11280
rect 25915 11172 26004 11200
rect 26436 11240 26608 11268
rect 25915 11169 25927 11172
rect 25869 11163 25927 11169
rect 24394 11132 24400 11144
rect 24136 11104 24400 11132
rect 24394 11092 24400 11104
rect 24452 11132 24458 11144
rect 24673 11135 24731 11141
rect 24673 11132 24685 11135
rect 24452 11104 24685 11132
rect 24452 11092 24458 11104
rect 24673 11101 24685 11104
rect 24719 11101 24731 11135
rect 24673 11095 24731 11101
rect 24765 11135 24823 11141
rect 24765 11101 24777 11135
rect 24811 11132 24823 11135
rect 24946 11132 24952 11144
rect 24811 11104 24952 11132
rect 24811 11101 24823 11104
rect 24765 11095 24823 11101
rect 24946 11092 24952 11104
rect 25004 11092 25010 11144
rect 25038 11092 25044 11144
rect 25096 11092 25102 11144
rect 25406 11092 25412 11144
rect 25464 11132 25470 11144
rect 25685 11135 25743 11141
rect 25685 11132 25697 11135
rect 25464 11104 25697 11132
rect 25464 11092 25470 11104
rect 25685 11101 25697 11104
rect 25731 11101 25743 11135
rect 25685 11095 25743 11101
rect 25777 11135 25835 11141
rect 25777 11101 25789 11135
rect 25823 11132 25835 11135
rect 26436 11132 26464 11240
rect 26602 11228 26608 11240
rect 26660 11228 26666 11280
rect 27338 11268 27344 11280
rect 26896 11240 27344 11268
rect 26510 11160 26516 11212
rect 26568 11160 26574 11212
rect 26896 11200 26924 11240
rect 27338 11228 27344 11240
rect 27396 11228 27402 11280
rect 29840 11268 29868 11296
rect 29012 11240 29868 11268
rect 29012 11209 29040 11240
rect 26620 11172 26924 11200
rect 26620 11132 26648 11172
rect 26896 11141 26924 11172
rect 27065 11203 27123 11209
rect 27065 11169 27077 11203
rect 27111 11200 27123 11203
rect 27157 11203 27215 11209
rect 27157 11200 27169 11203
rect 27111 11172 27169 11200
rect 27111 11169 27123 11172
rect 27065 11163 27123 11169
rect 27157 11169 27169 11172
rect 27203 11200 27215 11203
rect 28997 11203 29055 11209
rect 28997 11200 29009 11203
rect 27203 11172 28396 11200
rect 27203 11169 27215 11172
rect 27157 11163 27215 11169
rect 25823 11104 26464 11132
rect 26528 11104 26648 11132
rect 26881 11135 26939 11141
rect 25823 11101 25835 11104
rect 25777 11095 25835 11101
rect 23198 11024 23204 11076
rect 23256 11024 23262 11076
rect 23339 11067 23397 11073
rect 23339 11033 23351 11067
rect 23385 11064 23397 11067
rect 23385 11036 24716 11064
rect 23385 11033 23397 11036
rect 23339 11027 23397 11033
rect 24688 11008 24716 11036
rect 25314 11024 25320 11076
rect 25372 11064 25378 11076
rect 25590 11064 25596 11076
rect 25372 11036 25596 11064
rect 25372 11024 25378 11036
rect 25590 11024 25596 11036
rect 25648 11024 25654 11076
rect 25866 11024 25872 11076
rect 25924 11064 25930 11076
rect 26053 11067 26111 11073
rect 26053 11064 26065 11067
rect 25924 11036 26065 11064
rect 25924 11024 25930 11036
rect 26053 11033 26065 11036
rect 26099 11033 26111 11067
rect 26053 11027 26111 11033
rect 26269 11067 26327 11073
rect 26269 11033 26281 11067
rect 26315 11064 26327 11067
rect 26528 11064 26556 11104
rect 26881 11101 26893 11135
rect 26927 11101 26939 11135
rect 26881 11095 26939 11101
rect 26970 11092 26976 11144
rect 27028 11132 27034 11144
rect 27525 11135 27583 11141
rect 27525 11132 27537 11135
rect 27028 11104 27537 11132
rect 27028 11092 27034 11104
rect 27525 11101 27537 11104
rect 27571 11101 27583 11135
rect 27525 11095 27583 11101
rect 27614 11092 27620 11144
rect 27672 11092 27678 11144
rect 27798 11092 27804 11144
rect 27856 11132 27862 11144
rect 28368 11141 28396 11172
rect 28552 11172 29009 11200
rect 28552 11141 28580 11172
rect 28997 11169 29009 11172
rect 29043 11169 29055 11203
rect 29914 11200 29920 11212
rect 28997 11163 29055 11169
rect 29104 11172 29920 11200
rect 29104 11141 29132 11172
rect 29914 11160 29920 11172
rect 29972 11160 29978 11212
rect 28077 11135 28135 11141
rect 28077 11132 28089 11135
rect 27856 11104 28089 11132
rect 27856 11092 27862 11104
rect 28077 11101 28089 11104
rect 28123 11101 28135 11135
rect 28077 11095 28135 11101
rect 28353 11135 28411 11141
rect 28353 11101 28365 11135
rect 28399 11101 28411 11135
rect 28353 11095 28411 11101
rect 28537 11135 28595 11141
rect 28537 11101 28549 11135
rect 28583 11101 28595 11135
rect 28537 11095 28595 11101
rect 28813 11135 28871 11141
rect 28813 11101 28825 11135
rect 28859 11101 28871 11135
rect 28813 11095 28871 11101
rect 29089 11135 29147 11141
rect 29089 11101 29101 11135
rect 29135 11101 29147 11135
rect 29089 11095 29147 11101
rect 26315 11036 26556 11064
rect 26315 11033 26327 11036
rect 26269 11027 26327 11033
rect 27246 11024 27252 11076
rect 27304 11064 27310 11076
rect 28552 11064 28580 11095
rect 27304 11036 28580 11064
rect 28828 11064 28856 11095
rect 29546 11092 29552 11144
rect 29604 11092 29610 11144
rect 29638 11092 29644 11144
rect 29696 11092 29702 11144
rect 29730 11092 29736 11144
rect 29788 11132 29794 11144
rect 29825 11135 29883 11141
rect 29825 11132 29837 11135
rect 29788 11104 29837 11132
rect 29788 11092 29794 11104
rect 29825 11101 29837 11104
rect 29871 11101 29883 11135
rect 29825 11095 29883 11101
rect 29748 11064 29776 11092
rect 28828 11036 29776 11064
rect 27304 11024 27310 11036
rect 23474 10996 23480 11008
rect 23032 10968 23480 10996
rect 23474 10956 23480 10968
rect 23532 10956 23538 11008
rect 23934 10956 23940 11008
rect 23992 10996 23998 11008
rect 24397 10999 24455 11005
rect 24397 10996 24409 10999
rect 23992 10968 24409 10996
rect 23992 10956 23998 10968
rect 24397 10965 24409 10968
rect 24443 10965 24455 10999
rect 24397 10959 24455 10965
rect 24670 10956 24676 11008
rect 24728 10956 24734 11008
rect 24857 10999 24915 11005
rect 24857 10965 24869 10999
rect 24903 10996 24915 10999
rect 25332 10996 25360 11024
rect 24903 10968 25360 10996
rect 24903 10965 24915 10968
rect 24857 10959 24915 10965
rect 26418 10956 26424 11008
rect 26476 10956 26482 11008
rect 26694 10956 26700 11008
rect 26752 10956 26758 11008
rect 26789 10999 26847 11005
rect 26789 10965 26801 10999
rect 26835 10996 26847 10999
rect 26878 10996 26884 11008
rect 26835 10968 26884 10996
rect 26835 10965 26847 10968
rect 26789 10959 26847 10965
rect 26878 10956 26884 10968
rect 26936 10956 26942 11008
rect 27338 10956 27344 11008
rect 27396 10996 27402 11008
rect 28629 10999 28687 11005
rect 28629 10996 28641 10999
rect 27396 10968 28641 10996
rect 27396 10956 27402 10968
rect 28629 10965 28641 10968
rect 28675 10965 28687 10999
rect 28629 10959 28687 10965
rect 30006 10956 30012 11008
rect 30064 10956 30070 11008
rect 1104 10906 38824 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 35594 10906
rect 35646 10854 35658 10906
rect 35710 10854 35722 10906
rect 35774 10854 35786 10906
rect 35838 10854 35850 10906
rect 35902 10854 38824 10906
rect 1104 10832 38824 10854
rect 20990 10752 20996 10804
rect 21048 10792 21054 10804
rect 21269 10795 21327 10801
rect 21269 10792 21281 10795
rect 21048 10764 21281 10792
rect 21048 10752 21054 10764
rect 21269 10761 21281 10764
rect 21315 10761 21327 10795
rect 21269 10755 21327 10761
rect 21818 10752 21824 10804
rect 21876 10752 21882 10804
rect 22830 10792 22836 10804
rect 22112 10764 22836 10792
rect 20806 10616 20812 10668
rect 20864 10616 20870 10668
rect 21453 10659 21511 10665
rect 21453 10625 21465 10659
rect 21499 10656 21511 10659
rect 21836 10656 21864 10752
rect 22112 10733 22140 10764
rect 22830 10752 22836 10764
rect 22888 10752 22894 10804
rect 23566 10752 23572 10804
rect 23624 10752 23630 10804
rect 23750 10752 23756 10804
rect 23808 10752 23814 10804
rect 23842 10752 23848 10804
rect 23900 10792 23906 10804
rect 25222 10792 25228 10804
rect 23900 10764 25228 10792
rect 23900 10752 23906 10764
rect 25222 10752 25228 10764
rect 25280 10752 25286 10804
rect 26326 10752 26332 10804
rect 26384 10752 26390 10804
rect 26418 10752 26424 10804
rect 26476 10792 26482 10804
rect 26970 10792 26976 10804
rect 26476 10764 26976 10792
rect 26476 10752 26482 10764
rect 26970 10752 26976 10764
rect 27028 10752 27034 10804
rect 27338 10752 27344 10804
rect 27396 10752 27402 10804
rect 27617 10795 27675 10801
rect 27617 10761 27629 10795
rect 27663 10792 27675 10795
rect 27798 10792 27804 10804
rect 27663 10764 27804 10792
rect 27663 10761 27675 10764
rect 27617 10755 27675 10761
rect 27798 10752 27804 10764
rect 27856 10752 27862 10804
rect 27890 10752 27896 10804
rect 27948 10752 27954 10804
rect 29549 10795 29607 10801
rect 29549 10761 29561 10795
rect 29595 10792 29607 10795
rect 29638 10792 29644 10804
rect 29595 10764 29644 10792
rect 29595 10761 29607 10764
rect 29549 10755 29607 10761
rect 29638 10752 29644 10764
rect 29696 10752 29702 10804
rect 22097 10727 22155 10733
rect 22097 10693 22109 10727
rect 22143 10693 22155 10727
rect 23382 10724 23388 10736
rect 23322 10696 23388 10724
rect 22097 10687 22155 10693
rect 23382 10684 23388 10696
rect 23440 10684 23446 10736
rect 24044 10696 24900 10724
rect 21499 10628 21864 10656
rect 21499 10625 21511 10628
rect 21453 10619 21511 10625
rect 23934 10616 23940 10668
rect 23992 10616 23998 10668
rect 24044 10665 24072 10696
rect 24872 10668 24900 10696
rect 26234 10684 26240 10736
rect 26292 10684 26298 10736
rect 26344 10724 26372 10752
rect 26344 10696 27016 10724
rect 24029 10659 24087 10665
rect 24029 10625 24041 10659
rect 24075 10625 24087 10659
rect 24029 10619 24087 10625
rect 24305 10659 24363 10665
rect 24305 10625 24317 10659
rect 24351 10625 24363 10659
rect 24305 10619 24363 10625
rect 20824 10588 20852 10616
rect 21821 10591 21879 10597
rect 21821 10588 21833 10591
rect 20824 10560 21833 10588
rect 21821 10557 21833 10560
rect 21867 10557 21879 10591
rect 24320 10588 24348 10619
rect 24854 10616 24860 10668
rect 24912 10616 24918 10668
rect 25866 10616 25872 10668
rect 25924 10656 25930 10668
rect 26988 10665 27016 10696
rect 27246 10684 27252 10736
rect 27304 10724 27310 10736
rect 27458 10727 27516 10733
rect 27458 10724 27470 10727
rect 27304 10696 27470 10724
rect 27304 10684 27310 10696
rect 27458 10693 27470 10696
rect 27504 10693 27516 10727
rect 27908 10724 27936 10752
rect 28077 10727 28135 10733
rect 28077 10724 28089 10727
rect 27908 10696 28089 10724
rect 27458 10687 27516 10693
rect 28077 10693 28089 10696
rect 28123 10693 28135 10727
rect 28077 10687 28135 10693
rect 28810 10684 28816 10736
rect 28868 10684 28874 10736
rect 26329 10659 26387 10665
rect 26329 10656 26341 10659
rect 25924 10628 26341 10656
rect 25924 10616 25930 10628
rect 26329 10625 26341 10628
rect 26375 10625 26387 10659
rect 26329 10619 26387 10625
rect 26973 10659 27031 10665
rect 26973 10625 26985 10659
rect 27019 10625 27031 10659
rect 26973 10619 27031 10625
rect 25682 10588 25688 10600
rect 24320 10560 25688 10588
rect 21821 10551 21879 10557
rect 25682 10548 25688 10560
rect 25740 10548 25746 10600
rect 27249 10591 27307 10597
rect 27249 10588 27261 10591
rect 27172 10560 27261 10588
rect 24213 10523 24271 10529
rect 24213 10489 24225 10523
rect 24259 10520 24271 10523
rect 24670 10520 24676 10532
rect 24259 10492 24676 10520
rect 24259 10489 24271 10492
rect 24213 10483 24271 10489
rect 24670 10480 24676 10492
rect 24728 10480 24734 10532
rect 27172 10464 27200 10560
rect 27249 10557 27261 10560
rect 27295 10557 27307 10591
rect 27249 10551 27307 10557
rect 27614 10548 27620 10600
rect 27672 10588 27678 10600
rect 27801 10591 27859 10597
rect 27801 10588 27813 10591
rect 27672 10560 27813 10588
rect 27672 10548 27678 10560
rect 27801 10557 27813 10560
rect 27847 10557 27859 10591
rect 27801 10551 27859 10557
rect 22462 10412 22468 10464
rect 22520 10452 22526 10464
rect 24949 10455 25007 10461
rect 24949 10452 24961 10455
rect 22520 10424 24961 10452
rect 22520 10412 22526 10424
rect 24949 10421 24961 10424
rect 24995 10452 25007 10455
rect 25958 10452 25964 10464
rect 24995 10424 25964 10452
rect 24995 10421 25007 10424
rect 24949 10415 25007 10421
rect 25958 10412 25964 10424
rect 26016 10412 26022 10464
rect 26513 10455 26571 10461
rect 26513 10421 26525 10455
rect 26559 10452 26571 10455
rect 26694 10452 26700 10464
rect 26559 10424 26700 10452
rect 26559 10421 26571 10424
rect 26513 10415 26571 10421
rect 26694 10412 26700 10424
rect 26752 10452 26758 10464
rect 27154 10452 27160 10464
rect 26752 10424 27160 10452
rect 26752 10412 26758 10424
rect 27154 10412 27160 10424
rect 27212 10412 27218 10464
rect 1104 10362 38824 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38824 10362
rect 1104 10288 38824 10310
rect 20806 10208 20812 10260
rect 20864 10248 20870 10260
rect 21085 10251 21143 10257
rect 21085 10248 21097 10251
rect 20864 10220 21097 10248
rect 20864 10208 20870 10220
rect 21085 10217 21097 10220
rect 21131 10217 21143 10251
rect 21085 10211 21143 10217
rect 23474 10208 23480 10260
rect 23532 10208 23538 10260
rect 25130 10248 25136 10260
rect 25056 10220 25136 10248
rect 24394 10072 24400 10124
rect 24452 10072 24458 10124
rect 24486 10072 24492 10124
rect 24544 10072 24550 10124
rect 24578 10072 24584 10124
rect 24636 10072 24642 10124
rect 24765 10115 24823 10121
rect 24765 10081 24777 10115
rect 24811 10112 24823 10115
rect 24946 10112 24952 10124
rect 24811 10084 24952 10112
rect 24811 10081 24823 10084
rect 24765 10075 24823 10081
rect 23290 10004 23296 10056
rect 23348 10004 23354 10056
rect 23661 10047 23719 10053
rect 23661 10013 23673 10047
rect 23707 10044 23719 10047
rect 24412 10044 24440 10072
rect 24673 10047 24731 10053
rect 24673 10044 24685 10047
rect 23707 10016 24685 10044
rect 23707 10013 23719 10016
rect 23661 10007 23719 10013
rect 24673 10013 24685 10016
rect 24719 10013 24731 10047
rect 24673 10007 24731 10013
rect 22462 9936 22468 9988
rect 22520 9976 22526 9988
rect 22557 9979 22615 9985
rect 22557 9976 22569 9979
rect 22520 9948 22569 9976
rect 22520 9936 22526 9948
rect 22557 9945 22569 9948
rect 22603 9945 22615 9979
rect 22557 9939 22615 9945
rect 22922 9936 22928 9988
rect 22980 9976 22986 9988
rect 23845 9979 23903 9985
rect 23845 9976 23857 9979
rect 22980 9948 23857 9976
rect 22980 9936 22986 9948
rect 23845 9945 23857 9948
rect 23891 9976 23903 9979
rect 24780 9976 24808 10075
rect 24946 10072 24952 10084
rect 25004 10072 25010 10124
rect 25056 10044 25084 10220
rect 25130 10208 25136 10220
rect 25188 10208 25194 10260
rect 25498 10248 25504 10260
rect 25240 10220 25504 10248
rect 25130 10072 25136 10124
rect 25188 10112 25194 10124
rect 25240 10112 25268 10220
rect 25498 10208 25504 10220
rect 25556 10208 25562 10260
rect 27522 10208 27528 10260
rect 27580 10208 27586 10260
rect 25188 10084 25268 10112
rect 25593 10115 25651 10121
rect 25188 10072 25194 10084
rect 25593 10081 25605 10115
rect 25639 10112 25651 10115
rect 25639 10084 26280 10112
rect 25639 10081 25651 10084
rect 25593 10075 25651 10081
rect 26252 10056 26280 10084
rect 28460 10084 28994 10112
rect 25225 10047 25283 10053
rect 25225 10044 25237 10047
rect 25056 10016 25237 10044
rect 25225 10013 25237 10016
rect 25271 10013 25283 10047
rect 25225 10007 25283 10013
rect 25317 10047 25375 10053
rect 25317 10013 25329 10047
rect 25363 10013 25375 10047
rect 25317 10007 25375 10013
rect 23891 9948 24808 9976
rect 25332 9976 25360 10007
rect 25406 10004 25412 10056
rect 25464 10044 25470 10056
rect 25501 10047 25559 10053
rect 25501 10044 25513 10047
rect 25464 10016 25513 10044
rect 25464 10004 25470 10016
rect 25501 10013 25513 10016
rect 25547 10013 25559 10047
rect 25685 10047 25743 10053
rect 25685 10044 25697 10047
rect 25501 10007 25559 10013
rect 25608 10016 25697 10044
rect 25332 9948 25544 9976
rect 23891 9945 23903 9948
rect 23845 9939 23903 9945
rect 25516 9920 25544 9948
rect 25608 9920 25636 10016
rect 25685 10013 25697 10016
rect 25731 10013 25743 10047
rect 25685 10007 25743 10013
rect 25774 10004 25780 10056
rect 25832 10004 25838 10056
rect 25958 10004 25964 10056
rect 26016 10044 26022 10056
rect 26016 10016 26096 10044
rect 26016 10004 26022 10016
rect 26068 9985 26096 10016
rect 26234 10004 26240 10056
rect 26292 10004 26298 10056
rect 28074 10004 28080 10056
rect 28132 10004 28138 10056
rect 28460 10053 28488 10084
rect 28445 10047 28503 10053
rect 28445 10013 28457 10047
rect 28491 10013 28503 10047
rect 28966 10044 28994 10084
rect 29549 10047 29607 10053
rect 29549 10044 29561 10047
rect 28966 10016 29561 10044
rect 28445 10007 28503 10013
rect 29549 10013 29561 10016
rect 29595 10013 29607 10047
rect 29549 10007 29607 10013
rect 30006 10004 30012 10056
rect 30064 10004 30070 10056
rect 30098 10004 30104 10056
rect 30156 10004 30162 10056
rect 26053 9979 26111 9985
rect 26053 9945 26065 9979
rect 26099 9945 26111 9979
rect 26053 9939 26111 9945
rect 27246 9936 27252 9988
rect 27304 9976 27310 9988
rect 27304 9948 28028 9976
rect 27304 9936 27310 9948
rect 22738 9868 22744 9920
rect 22796 9868 22802 9920
rect 24946 9868 24952 9920
rect 25004 9868 25010 9920
rect 25498 9868 25504 9920
rect 25556 9868 25562 9920
rect 25590 9868 25596 9920
rect 25648 9868 25654 9920
rect 25958 9868 25964 9920
rect 26016 9868 26022 9920
rect 27706 9868 27712 9920
rect 27764 9908 27770 9920
rect 27893 9911 27951 9917
rect 27893 9908 27905 9911
rect 27764 9880 27905 9908
rect 27764 9868 27770 9880
rect 27893 9877 27905 9880
rect 27939 9877 27951 9911
rect 28000 9908 28028 9948
rect 28166 9936 28172 9988
rect 28224 9936 28230 9988
rect 28261 9979 28319 9985
rect 28261 9945 28273 9979
rect 28307 9976 28319 9979
rect 28626 9976 28632 9988
rect 28307 9948 28632 9976
rect 28307 9945 28319 9948
rect 28261 9939 28319 9945
rect 28626 9936 28632 9948
rect 28684 9936 28690 9988
rect 28718 9936 28724 9988
rect 28776 9936 28782 9988
rect 28905 9979 28963 9985
rect 28905 9945 28917 9979
rect 28951 9976 28963 9979
rect 30024 9976 30052 10004
rect 28951 9948 30052 9976
rect 28951 9945 28963 9948
rect 28905 9939 28963 9945
rect 28537 9911 28595 9917
rect 28537 9908 28549 9911
rect 28000 9880 28549 9908
rect 27893 9871 27951 9877
rect 28537 9877 28549 9880
rect 28583 9877 28595 9911
rect 28537 9871 28595 9877
rect 1104 9818 38824 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 35594 9818
rect 35646 9766 35658 9818
rect 35710 9766 35722 9818
rect 35774 9766 35786 9818
rect 35838 9766 35850 9818
rect 35902 9766 38824 9818
rect 1104 9744 38824 9766
rect 22940 9676 23980 9704
rect 22940 9636 22968 9676
rect 22296 9608 22968 9636
rect 22296 9577 22324 9608
rect 23014 9596 23020 9648
rect 23072 9636 23078 9648
rect 23952 9636 23980 9676
rect 24946 9664 24952 9716
rect 25004 9704 25010 9716
rect 25004 9676 25636 9704
rect 25004 9664 25010 9676
rect 24578 9636 24584 9648
rect 23072 9608 23138 9636
rect 23952 9608 24584 9636
rect 23072 9596 23078 9608
rect 24578 9596 24584 9608
rect 24636 9596 24642 9648
rect 25038 9596 25044 9648
rect 25096 9636 25102 9648
rect 25096 9608 25344 9636
rect 25096 9596 25102 9608
rect 25271 9605 25344 9608
rect 22281 9571 22339 9577
rect 22281 9537 22293 9571
rect 22327 9537 22339 9571
rect 22281 9531 22339 9537
rect 22465 9571 22523 9577
rect 22465 9537 22477 9571
rect 22511 9568 22523 9571
rect 22738 9568 22744 9580
rect 22511 9540 22744 9568
rect 22511 9537 22523 9540
rect 22465 9531 22523 9537
rect 22738 9528 22744 9540
rect 22796 9528 22802 9580
rect 24596 9568 24624 9596
rect 24857 9571 24915 9577
rect 24857 9568 24869 9571
rect 24596 9540 24869 9568
rect 24857 9537 24869 9540
rect 24903 9537 24915 9571
rect 25271 9571 25283 9605
rect 25317 9571 25344 9605
rect 25498 9596 25504 9648
rect 25556 9596 25562 9648
rect 25608 9636 25636 9676
rect 25682 9664 25688 9716
rect 25740 9664 25746 9716
rect 25866 9664 25872 9716
rect 25924 9664 25930 9716
rect 26142 9704 26148 9716
rect 26068 9676 26148 9704
rect 26068 9636 26096 9676
rect 26142 9664 26148 9676
rect 26200 9664 26206 9716
rect 26234 9664 26240 9716
rect 26292 9704 26298 9716
rect 29181 9707 29239 9713
rect 29181 9704 29193 9707
rect 26292 9676 29193 9704
rect 26292 9664 26298 9676
rect 29181 9673 29193 9676
rect 29227 9704 29239 9707
rect 30098 9704 30104 9716
rect 29227 9676 30104 9704
rect 29227 9673 29239 9676
rect 29181 9667 29239 9673
rect 30098 9664 30104 9676
rect 30156 9664 30162 9716
rect 25608 9608 26096 9636
rect 25792 9577 25820 9608
rect 25271 9565 25344 9571
rect 24857 9531 24915 9537
rect 24302 9460 24308 9512
rect 24360 9460 24366 9512
rect 24581 9503 24639 9509
rect 24581 9469 24593 9503
rect 24627 9469 24639 9503
rect 24581 9463 24639 9469
rect 24596 9432 24624 9463
rect 24670 9460 24676 9512
rect 24728 9500 24734 9512
rect 25041 9503 25099 9509
rect 25041 9500 25053 9503
rect 24728 9472 25053 9500
rect 24728 9460 24734 9472
rect 25041 9469 25053 9472
rect 25087 9469 25099 9503
rect 25316 9500 25344 9565
rect 25777 9571 25835 9577
rect 25777 9537 25789 9571
rect 25823 9537 25835 9571
rect 25777 9531 25835 9537
rect 25866 9528 25872 9580
rect 25924 9568 25930 9580
rect 26053 9571 26111 9577
rect 26053 9568 26065 9571
rect 25924 9540 26065 9568
rect 25924 9528 25930 9540
rect 26053 9537 26065 9540
rect 26099 9537 26111 9571
rect 26053 9531 26111 9537
rect 26142 9528 26148 9580
rect 26200 9528 26206 9580
rect 26252 9577 26280 9664
rect 27246 9636 27252 9648
rect 26528 9608 27252 9636
rect 26528 9577 26556 9608
rect 26237 9571 26295 9577
rect 26237 9537 26249 9571
rect 26283 9537 26295 9571
rect 26237 9531 26295 9537
rect 26421 9571 26479 9577
rect 26421 9537 26433 9571
rect 26467 9537 26479 9571
rect 26421 9531 26479 9537
rect 26513 9571 26571 9577
rect 26513 9537 26525 9571
rect 26559 9537 26571 9571
rect 26513 9531 26571 9537
rect 25958 9500 25964 9512
rect 25316 9472 25964 9500
rect 25041 9463 25099 9469
rect 25958 9460 25964 9472
rect 26016 9460 26022 9512
rect 25498 9432 25504 9444
rect 24596 9404 25504 9432
rect 25498 9392 25504 9404
rect 25556 9392 25562 9444
rect 21726 9324 21732 9376
rect 21784 9364 21790 9376
rect 22097 9367 22155 9373
rect 22097 9364 22109 9367
rect 21784 9336 22109 9364
rect 21784 9324 21790 9336
rect 22097 9333 22109 9336
rect 22143 9333 22155 9367
rect 22097 9327 22155 9333
rect 22830 9324 22836 9376
rect 22888 9324 22894 9376
rect 24670 9324 24676 9376
rect 24728 9324 24734 9376
rect 25133 9367 25191 9373
rect 25133 9333 25145 9367
rect 25179 9364 25191 9367
rect 25222 9364 25228 9376
rect 25179 9336 25228 9364
rect 25179 9333 25191 9336
rect 25133 9327 25191 9333
rect 25222 9324 25228 9336
rect 25280 9324 25286 9376
rect 25314 9324 25320 9376
rect 25372 9324 25378 9376
rect 25406 9324 25412 9376
rect 25464 9364 25470 9376
rect 26436 9364 26464 9531
rect 26602 9528 26608 9580
rect 26660 9528 26666 9580
rect 26804 9577 26832 9608
rect 27246 9596 27252 9608
rect 27304 9596 27310 9648
rect 27706 9596 27712 9648
rect 27764 9596 27770 9648
rect 28258 9596 28264 9648
rect 28316 9596 28322 9648
rect 26789 9571 26847 9577
rect 26789 9537 26801 9571
rect 26835 9537 26847 9571
rect 26789 9531 26847 9537
rect 26973 9571 27031 9577
rect 26973 9537 26985 9571
rect 27019 9537 27031 9571
rect 26973 9531 27031 9537
rect 26694 9460 26700 9512
rect 26752 9460 26758 9512
rect 26878 9460 26884 9512
rect 26936 9500 26942 9512
rect 26988 9500 27016 9531
rect 26936 9472 27016 9500
rect 26936 9460 26942 9472
rect 27062 9460 27068 9512
rect 27120 9460 27126 9512
rect 27430 9500 27436 9512
rect 27264 9472 27436 9500
rect 26712 9432 26740 9460
rect 27264 9432 27292 9472
rect 27430 9460 27436 9472
rect 27488 9460 27494 9512
rect 26712 9404 27292 9432
rect 27338 9392 27344 9444
rect 27396 9392 27402 9444
rect 25464 9336 26464 9364
rect 25464 9324 25470 9336
rect 26510 9324 26516 9376
rect 26568 9364 26574 9376
rect 26789 9367 26847 9373
rect 26789 9364 26801 9367
rect 26568 9336 26801 9364
rect 26568 9324 26574 9336
rect 26789 9333 26801 9336
rect 26835 9364 26847 9367
rect 26970 9364 26976 9376
rect 26835 9336 26976 9364
rect 26835 9333 26847 9336
rect 26789 9327 26847 9333
rect 26970 9324 26976 9336
rect 27028 9324 27034 9376
rect 27154 9324 27160 9376
rect 27212 9364 27218 9376
rect 28442 9364 28448 9376
rect 27212 9336 28448 9364
rect 27212 9324 27218 9336
rect 28442 9324 28448 9336
rect 28500 9324 28506 9376
rect 1104 9274 38824 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38824 9274
rect 1104 9200 38824 9222
rect 22925 9163 22983 9169
rect 22925 9129 22937 9163
rect 22971 9160 22983 9163
rect 23290 9160 23296 9172
rect 22971 9132 23296 9160
rect 22971 9129 22983 9132
rect 22925 9123 22983 9129
rect 23290 9120 23296 9132
rect 23348 9120 23354 9172
rect 24121 9163 24179 9169
rect 24121 9129 24133 9163
rect 24167 9160 24179 9163
rect 24302 9160 24308 9172
rect 24167 9132 24308 9160
rect 24167 9129 24179 9132
rect 24121 9123 24179 9129
rect 24302 9120 24308 9132
rect 24360 9120 24366 9172
rect 24578 9120 24584 9172
rect 24636 9120 24642 9172
rect 24670 9120 24676 9172
rect 24728 9120 24734 9172
rect 25774 9120 25780 9172
rect 25832 9160 25838 9172
rect 26786 9160 26792 9172
rect 25832 9132 26792 9160
rect 25832 9120 25838 9132
rect 26786 9120 26792 9132
rect 26844 9120 26850 9172
rect 28258 9160 28264 9172
rect 27908 9132 28264 9160
rect 23845 9095 23903 9101
rect 23845 9061 23857 9095
rect 23891 9092 23903 9095
rect 24596 9092 24624 9120
rect 23891 9064 24624 9092
rect 23891 9061 23903 9064
rect 23845 9055 23903 9061
rect 21177 9027 21235 9033
rect 21177 8993 21189 9027
rect 21223 9024 21235 9027
rect 21818 9024 21824 9036
rect 21223 8996 21824 9024
rect 21223 8993 21235 8996
rect 21177 8987 21235 8993
rect 21818 8984 21824 8996
rect 21876 8984 21882 9036
rect 22830 8984 22836 9036
rect 22888 9024 22894 9036
rect 23014 9024 23020 9036
rect 22888 8996 23020 9024
rect 22888 8984 22894 8996
rect 23014 8984 23020 8996
rect 23072 9024 23078 9036
rect 23201 9027 23259 9033
rect 23201 9024 23213 9027
rect 23072 8996 23213 9024
rect 23072 8984 23078 8996
rect 23201 8993 23213 8996
rect 23247 8993 23259 9027
rect 23201 8987 23259 8993
rect 22554 8916 22560 8968
rect 22612 8956 22618 8968
rect 22922 8956 22928 8968
rect 22612 8928 22928 8956
rect 22612 8916 22618 8928
rect 22922 8916 22928 8928
rect 22980 8916 22986 8968
rect 23937 8959 23995 8965
rect 23937 8925 23949 8959
rect 23983 8956 23995 8959
rect 24688 8956 24716 9120
rect 26694 9092 26700 9104
rect 26160 9064 26700 9092
rect 25498 8984 25504 9036
rect 25556 9024 25562 9036
rect 26160 9033 26188 9064
rect 26694 9052 26700 9064
rect 26752 9052 26758 9104
rect 26804 9092 26832 9120
rect 27908 9092 27936 9132
rect 28258 9120 28264 9132
rect 28316 9120 28322 9172
rect 28534 9120 28540 9172
rect 28592 9120 28598 9172
rect 28626 9120 28632 9172
rect 28684 9160 28690 9172
rect 29825 9163 29883 9169
rect 29825 9160 29837 9163
rect 28684 9132 29837 9160
rect 28684 9120 28690 9132
rect 29825 9129 29837 9132
rect 29871 9129 29883 9163
rect 29825 9123 29883 9129
rect 30006 9120 30012 9172
rect 30064 9120 30070 9172
rect 28644 9092 28672 9120
rect 26804 9064 27936 9092
rect 28000 9064 28672 9092
rect 29549 9095 29607 9101
rect 26145 9027 26203 9033
rect 26145 9024 26157 9027
rect 25556 8996 26157 9024
rect 25556 8984 25562 8996
rect 26145 8993 26157 8996
rect 26191 8993 26203 9027
rect 26881 9027 26939 9033
rect 26145 8987 26203 8993
rect 26252 8996 26464 9024
rect 23983 8928 24716 8956
rect 23983 8925 23995 8928
rect 23937 8919 23995 8925
rect 21450 8848 21456 8900
rect 21508 8848 21514 8900
rect 25774 8888 25780 8900
rect 25438 8860 25780 8888
rect 25774 8848 25780 8860
rect 25832 8848 25838 8900
rect 25869 8891 25927 8897
rect 25869 8857 25881 8891
rect 25915 8888 25927 8891
rect 26252 8888 26280 8996
rect 26329 8959 26387 8965
rect 26329 8925 26341 8959
rect 26375 8925 26387 8959
rect 26436 8956 26464 8996
rect 26881 8993 26893 9027
rect 26927 9024 26939 9027
rect 27249 9027 27307 9033
rect 27249 9024 27261 9027
rect 26927 8996 27261 9024
rect 26927 8993 26939 8996
rect 26881 8987 26939 8993
rect 27249 8993 27261 8996
rect 27295 8993 27307 9027
rect 27249 8987 27307 8993
rect 27338 8984 27344 9036
rect 27396 9024 27402 9036
rect 27617 9027 27675 9033
rect 27617 9024 27629 9027
rect 27396 8996 27629 9024
rect 27396 8984 27402 8996
rect 27617 8993 27629 8996
rect 27663 8993 27675 9027
rect 27617 8987 27675 8993
rect 26973 8959 27031 8965
rect 26973 8956 26985 8959
rect 26436 8928 26985 8956
rect 26329 8919 26387 8925
rect 26973 8925 26985 8928
rect 27019 8925 27031 8959
rect 26973 8919 27031 8925
rect 27157 8959 27215 8965
rect 27157 8925 27169 8959
rect 27203 8956 27215 8959
rect 28000 8956 28028 9064
rect 29549 9061 29561 9095
rect 29595 9092 29607 9095
rect 29730 9092 29736 9104
rect 29595 9064 29736 9092
rect 29595 9061 29607 9064
rect 29549 9055 29607 9061
rect 29730 9052 29736 9064
rect 29788 9092 29794 9104
rect 30024 9092 30052 9120
rect 29788 9064 30052 9092
rect 29788 9052 29794 9064
rect 28074 8984 28080 9036
rect 28132 9024 28138 9036
rect 28261 9027 28319 9033
rect 28261 9024 28273 9027
rect 28132 8996 28273 9024
rect 28132 8984 28138 8996
rect 28261 8993 28273 8996
rect 28307 9024 28319 9027
rect 28307 8996 29868 9024
rect 28307 8993 28319 8996
rect 28261 8987 28319 8993
rect 27203 8928 28028 8956
rect 27203 8925 27215 8928
rect 27157 8919 27215 8925
rect 25915 8860 26280 8888
rect 25915 8857 25927 8860
rect 25869 8851 25927 8857
rect 24397 8823 24455 8829
rect 24397 8789 24409 8823
rect 24443 8820 24455 8823
rect 25590 8820 25596 8832
rect 24443 8792 25596 8820
rect 24443 8789 24455 8792
rect 24397 8783 24455 8789
rect 25590 8780 25596 8792
rect 25648 8820 25654 8832
rect 26142 8820 26148 8832
rect 25648 8792 26148 8820
rect 25648 8780 25654 8792
rect 26142 8780 26148 8792
rect 26200 8820 26206 8832
rect 26344 8820 26372 8919
rect 28166 8916 28172 8968
rect 28224 8956 28230 8968
rect 29840 8965 29868 8996
rect 28353 8959 28411 8965
rect 28353 8956 28365 8959
rect 28224 8928 28365 8956
rect 28224 8916 28230 8928
rect 28353 8925 28365 8928
rect 28399 8925 28411 8959
rect 28353 8919 28411 8925
rect 28629 8959 28687 8965
rect 28629 8925 28641 8959
rect 28675 8925 28687 8959
rect 28629 8919 28687 8925
rect 29825 8959 29883 8965
rect 29825 8925 29837 8959
rect 29871 8925 29883 8959
rect 29825 8919 29883 8925
rect 30009 8959 30067 8965
rect 30009 8925 30021 8959
rect 30055 8925 30067 8959
rect 30009 8919 30067 8925
rect 27709 8891 27767 8897
rect 27709 8857 27721 8891
rect 27755 8857 27767 8891
rect 27985 8891 28043 8897
rect 27985 8888 27997 8891
rect 27709 8851 27767 8857
rect 27816 8860 27997 8888
rect 27062 8820 27068 8832
rect 26200 8792 27068 8820
rect 26200 8780 26206 8792
rect 27062 8780 27068 8792
rect 27120 8820 27126 8832
rect 27724 8820 27752 8851
rect 27816 8832 27844 8860
rect 27985 8857 27997 8860
rect 28031 8888 28043 8891
rect 28644 8888 28672 8919
rect 28031 8860 28672 8888
rect 28031 8857 28043 8860
rect 27985 8851 28043 8857
rect 28718 8848 28724 8900
rect 28776 8888 28782 8900
rect 30024 8888 30052 8919
rect 28776 8860 30052 8888
rect 28776 8848 28782 8860
rect 27120 8792 27752 8820
rect 27120 8780 27126 8792
rect 27798 8780 27804 8832
rect 27856 8780 27862 8832
rect 27890 8780 27896 8832
rect 27948 8780 27954 8832
rect 28074 8780 28080 8832
rect 28132 8780 28138 8832
rect 28905 8823 28963 8829
rect 28905 8789 28917 8823
rect 28951 8820 28963 8823
rect 29546 8820 29552 8832
rect 28951 8792 29552 8820
rect 28951 8789 28963 8792
rect 28905 8783 28963 8789
rect 29546 8780 29552 8792
rect 29604 8780 29610 8832
rect 1104 8730 38824 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 35594 8730
rect 35646 8678 35658 8730
rect 35710 8678 35722 8730
rect 35774 8678 35786 8730
rect 35838 8678 35850 8730
rect 35902 8678 38824 8730
rect 1104 8656 38824 8678
rect 21450 8576 21456 8628
rect 21508 8576 21514 8628
rect 21726 8576 21732 8628
rect 21784 8576 21790 8628
rect 25869 8619 25927 8625
rect 21836 8588 24164 8616
rect 21637 8483 21695 8489
rect 21637 8449 21649 8483
rect 21683 8480 21695 8483
rect 21744 8480 21772 8576
rect 21836 8492 21864 8588
rect 22554 8508 22560 8560
rect 22612 8508 22618 8560
rect 21683 8452 21772 8480
rect 21683 8449 21695 8452
rect 21637 8443 21695 8449
rect 21818 8440 21824 8492
rect 21876 8440 21882 8492
rect 24136 8489 24164 8588
rect 25869 8585 25881 8619
rect 25915 8616 25927 8619
rect 25915 8588 27384 8616
rect 25915 8585 25927 8588
rect 25869 8579 25927 8585
rect 25774 8548 25780 8560
rect 25622 8520 25780 8548
rect 25774 8508 25780 8520
rect 25832 8508 25838 8560
rect 26237 8551 26295 8557
rect 26237 8517 26249 8551
rect 26283 8548 26295 8551
rect 27356 8548 27384 8588
rect 27430 8576 27436 8628
rect 27488 8616 27494 8628
rect 28902 8616 28908 8628
rect 27488 8588 28908 8616
rect 27488 8576 27494 8588
rect 28902 8576 28908 8588
rect 28960 8616 28966 8628
rect 28960 8588 29960 8616
rect 28960 8576 28966 8588
rect 27890 8548 27896 8560
rect 26283 8520 27200 8548
rect 27356 8520 27896 8548
rect 26283 8517 26295 8520
rect 26237 8511 26295 8517
rect 23845 8483 23903 8489
rect 23845 8449 23857 8483
rect 23891 8449 23903 8483
rect 23845 8443 23903 8449
rect 24121 8483 24179 8489
rect 24121 8449 24133 8483
rect 24167 8449 24179 8483
rect 24121 8443 24179 8449
rect 26145 8483 26203 8489
rect 26145 8449 26157 8483
rect 26191 8449 26203 8483
rect 26145 8443 26203 8449
rect 22094 8372 22100 8424
rect 22152 8372 22158 8424
rect 23566 8236 23572 8288
rect 23624 8236 23630 8288
rect 23658 8236 23664 8288
rect 23716 8236 23722 8288
rect 23860 8276 23888 8443
rect 24026 8372 24032 8424
rect 24084 8372 24090 8424
rect 24397 8415 24455 8421
rect 24397 8381 24409 8415
rect 24443 8412 24455 8415
rect 25961 8415 26019 8421
rect 25961 8412 25973 8415
rect 24443 8384 25973 8412
rect 24443 8381 24455 8384
rect 24397 8375 24455 8381
rect 25961 8381 25973 8384
rect 26007 8381 26019 8415
rect 26160 8412 26188 8443
rect 26326 8440 26332 8492
rect 26384 8440 26390 8492
rect 26418 8440 26424 8492
rect 26476 8489 26482 8492
rect 26476 8483 26505 8489
rect 26493 8449 26505 8483
rect 27172 8480 27200 8520
rect 27632 8492 27660 8520
rect 27890 8508 27896 8520
rect 27948 8508 27954 8560
rect 28258 8508 28264 8560
rect 28316 8548 28322 8560
rect 28316 8520 28474 8548
rect 28316 8508 28322 8520
rect 29638 8508 29644 8560
rect 29696 8508 29702 8560
rect 27522 8480 27528 8492
rect 27172 8452 27528 8480
rect 26476 8443 26505 8449
rect 26476 8440 26482 8443
rect 27522 8440 27528 8452
rect 27580 8440 27586 8492
rect 27614 8440 27620 8492
rect 27672 8480 27678 8492
rect 27709 8483 27767 8489
rect 27709 8480 27721 8483
rect 27672 8452 27721 8480
rect 27672 8440 27678 8452
rect 27709 8449 27721 8452
rect 27755 8449 27767 8483
rect 27709 8443 27767 8449
rect 27798 8440 27804 8492
rect 27856 8440 27862 8492
rect 27985 8483 28043 8489
rect 27985 8449 27997 8483
rect 28031 8480 28043 8483
rect 28074 8480 28080 8492
rect 28031 8452 28080 8480
rect 28031 8449 28043 8452
rect 27985 8443 28043 8449
rect 28074 8440 28080 8452
rect 28132 8480 28138 8492
rect 29932 8489 29960 8588
rect 38194 8576 38200 8628
rect 38252 8616 38258 8628
rect 38289 8619 38347 8625
rect 38289 8616 38301 8619
rect 38252 8588 38301 8616
rect 38252 8576 38258 8588
rect 38289 8585 38301 8588
rect 38335 8585 38347 8619
rect 38289 8579 38347 8585
rect 30377 8551 30435 8557
rect 30377 8548 30389 8551
rect 30024 8520 30389 8548
rect 30024 8492 30052 8520
rect 30377 8517 30389 8520
rect 30423 8517 30435 8551
rect 30377 8511 30435 8517
rect 29917 8483 29975 8489
rect 28132 8452 28488 8480
rect 28132 8440 28138 8452
rect 26605 8415 26663 8421
rect 26160 8384 26556 8412
rect 25961 8375 26019 8381
rect 26528 8344 26556 8384
rect 26605 8381 26617 8415
rect 26651 8412 26663 8415
rect 26973 8415 27031 8421
rect 26973 8412 26985 8415
rect 26651 8384 26985 8412
rect 26651 8381 26663 8384
rect 26605 8375 26663 8381
rect 26973 8381 26985 8384
rect 27019 8381 27031 8415
rect 27816 8412 27844 8440
rect 27816 8384 28212 8412
rect 26973 8375 27031 8381
rect 26878 8344 26884 8356
rect 26528 8316 26884 8344
rect 26878 8304 26884 8316
rect 26936 8344 26942 8356
rect 27709 8347 27767 8353
rect 27709 8344 27721 8347
rect 26936 8316 27721 8344
rect 26936 8304 26942 8316
rect 27709 8313 27721 8316
rect 27755 8313 27767 8347
rect 27709 8307 27767 8313
rect 24486 8276 24492 8288
rect 23860 8248 24492 8276
rect 24486 8236 24492 8248
rect 24544 8236 24550 8288
rect 28184 8285 28212 8384
rect 28460 8288 28488 8452
rect 29917 8449 29929 8483
rect 29963 8449 29975 8483
rect 29917 8443 29975 8449
rect 30006 8440 30012 8492
rect 30064 8440 30070 8492
rect 30190 8440 30196 8492
rect 30248 8440 30254 8492
rect 30285 8483 30343 8489
rect 30285 8449 30297 8483
rect 30331 8449 30343 8483
rect 30285 8443 30343 8449
rect 28626 8372 28632 8424
rect 28684 8412 28690 8424
rect 30300 8412 30328 8443
rect 30558 8440 30564 8492
rect 30616 8440 30622 8492
rect 38381 8483 38439 8489
rect 38381 8449 38393 8483
rect 38427 8480 38439 8483
rect 38427 8452 38884 8480
rect 38427 8449 38439 8452
rect 38381 8443 38439 8449
rect 28684 8384 30328 8412
rect 28684 8372 28690 8384
rect 38856 8356 38884 8452
rect 38838 8304 38844 8356
rect 38896 8304 38902 8356
rect 28169 8279 28227 8285
rect 28169 8245 28181 8279
rect 28215 8276 28227 8279
rect 28350 8276 28356 8288
rect 28215 8248 28356 8276
rect 28215 8245 28227 8248
rect 28169 8239 28227 8245
rect 28350 8236 28356 8248
rect 28408 8236 28414 8288
rect 28442 8236 28448 8288
rect 28500 8236 28506 8288
rect 29822 8236 29828 8288
rect 29880 8276 29886 8288
rect 30009 8279 30067 8285
rect 30009 8276 30021 8279
rect 29880 8248 30021 8276
rect 29880 8236 29886 8248
rect 30009 8245 30021 8248
rect 30055 8245 30067 8279
rect 30009 8239 30067 8245
rect 1104 8186 38824 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38824 8186
rect 1104 8112 38824 8134
rect 20806 8032 20812 8084
rect 20864 8072 20870 8084
rect 21269 8075 21327 8081
rect 21269 8072 21281 8075
rect 20864 8044 21281 8072
rect 20864 8032 20870 8044
rect 21269 8041 21281 8044
rect 21315 8072 21327 8075
rect 21818 8072 21824 8084
rect 21315 8044 21824 8072
rect 21315 8041 21327 8044
rect 21269 8035 21327 8041
rect 21818 8032 21824 8044
rect 21876 8032 21882 8084
rect 22094 8032 22100 8084
rect 22152 8072 22158 8084
rect 22649 8075 22707 8081
rect 22649 8072 22661 8075
rect 22152 8044 22661 8072
rect 22152 8032 22158 8044
rect 22649 8041 22661 8044
rect 22695 8041 22707 8075
rect 22649 8035 22707 8041
rect 23201 8075 23259 8081
rect 23201 8041 23213 8075
rect 23247 8072 23259 8075
rect 23290 8072 23296 8084
rect 23247 8044 23296 8072
rect 23247 8041 23259 8044
rect 23201 8035 23259 8041
rect 23290 8032 23296 8044
rect 23348 8032 23354 8084
rect 23658 8032 23664 8084
rect 23716 8032 23722 8084
rect 24026 8032 24032 8084
rect 24084 8072 24090 8084
rect 24121 8075 24179 8081
rect 24121 8072 24133 8075
rect 24084 8044 24133 8072
rect 24084 8032 24090 8044
rect 24121 8041 24133 8044
rect 24167 8041 24179 8075
rect 24121 8035 24179 8041
rect 27062 8032 27068 8084
rect 27120 8072 27126 8084
rect 27341 8075 27399 8081
rect 27341 8072 27353 8075
rect 27120 8044 27353 8072
rect 27120 8032 27126 8044
rect 27341 8041 27353 8044
rect 27387 8072 27399 8075
rect 27430 8072 27436 8084
rect 27387 8044 27436 8072
rect 27387 8041 27399 8044
rect 27341 8035 27399 8041
rect 27430 8032 27436 8044
rect 27488 8032 27494 8084
rect 27982 8032 27988 8084
rect 28040 8072 28046 8084
rect 28258 8072 28264 8084
rect 28040 8044 28264 8072
rect 28040 8032 28046 8044
rect 28258 8032 28264 8044
rect 28316 8072 28322 8084
rect 29270 8072 29276 8084
rect 28316 8044 29276 8072
rect 28316 8032 28322 8044
rect 29270 8032 29276 8044
rect 29328 8032 29334 8084
rect 29638 8032 29644 8084
rect 29696 8072 29702 8084
rect 30193 8075 30251 8081
rect 30193 8072 30205 8075
rect 29696 8044 30205 8072
rect 29696 8032 29702 8044
rect 30193 8041 30205 8044
rect 30239 8041 30251 8075
rect 30193 8035 30251 8041
rect 30558 8032 30564 8084
rect 30616 8072 30622 8084
rect 30929 8075 30987 8081
rect 30929 8072 30941 8075
rect 30616 8044 30941 8072
rect 30616 8032 30622 8044
rect 30929 8041 30941 8044
rect 30975 8041 30987 8075
rect 30929 8035 30987 8041
rect 23676 8004 23704 8032
rect 22848 7976 23704 8004
rect 25976 7976 29776 8004
rect 22462 7828 22468 7880
rect 22520 7868 22526 7880
rect 22848 7877 22876 7976
rect 23109 7939 23167 7945
rect 23109 7905 23121 7939
rect 23155 7936 23167 7939
rect 23566 7936 23572 7948
rect 23155 7908 23572 7936
rect 23155 7905 23167 7908
rect 23109 7899 23167 7905
rect 23566 7896 23572 7908
rect 23624 7896 23630 7948
rect 22557 7871 22615 7877
rect 22557 7868 22569 7871
rect 22520 7840 22569 7868
rect 22520 7828 22526 7840
rect 22557 7837 22569 7840
rect 22603 7837 22615 7871
rect 22557 7831 22615 7837
rect 22833 7871 22891 7877
rect 22833 7837 22845 7871
rect 22879 7837 22891 7871
rect 22833 7831 22891 7837
rect 23014 7828 23020 7880
rect 23072 7868 23078 7880
rect 25976 7877 26004 7976
rect 29748 7948 29776 7976
rect 27798 7896 27804 7948
rect 27856 7936 27862 7948
rect 28626 7936 28632 7948
rect 27856 7908 28632 7936
rect 27856 7896 27862 7908
rect 23201 7871 23259 7877
rect 23201 7868 23213 7871
rect 23072 7840 23213 7868
rect 23072 7828 23078 7840
rect 23201 7837 23213 7840
rect 23247 7837 23259 7871
rect 23201 7831 23259 7837
rect 25961 7871 26019 7877
rect 25961 7837 25973 7871
rect 26007 7837 26019 7871
rect 25961 7831 26019 7837
rect 26050 7828 26056 7880
rect 26108 7828 26114 7880
rect 28092 7877 28120 7908
rect 28626 7896 28632 7908
rect 28684 7896 28690 7948
rect 29546 7896 29552 7948
rect 29604 7896 29610 7948
rect 29730 7896 29736 7948
rect 29788 7896 29794 7948
rect 27985 7871 28043 7877
rect 27985 7837 27997 7871
rect 28031 7837 28043 7871
rect 27985 7831 28043 7837
rect 28077 7871 28135 7877
rect 28077 7837 28089 7871
rect 28123 7837 28135 7871
rect 28077 7831 28135 7837
rect 22922 7760 22928 7812
rect 22980 7760 22986 7812
rect 24486 7760 24492 7812
rect 24544 7800 24550 7812
rect 24544 7772 25820 7800
rect 24544 7760 24550 7772
rect 23385 7735 23443 7741
rect 23385 7701 23397 7735
rect 23431 7732 23443 7735
rect 25406 7732 25412 7744
rect 23431 7704 25412 7732
rect 23431 7701 23443 7704
rect 23385 7695 23443 7701
rect 25406 7692 25412 7704
rect 25464 7692 25470 7744
rect 25792 7741 25820 7772
rect 27890 7760 27896 7812
rect 27948 7800 27954 7812
rect 28000 7800 28028 7831
rect 28350 7828 28356 7880
rect 28408 7828 28414 7880
rect 28997 7871 29055 7877
rect 28997 7837 29009 7871
rect 29043 7868 29055 7871
rect 29917 7871 29975 7877
rect 29917 7868 29929 7871
rect 29043 7840 29929 7868
rect 29043 7837 29055 7840
rect 28997 7831 29055 7837
rect 29917 7837 29929 7840
rect 29963 7837 29975 7871
rect 29917 7831 29975 7837
rect 30006 7828 30012 7880
rect 30064 7828 30070 7880
rect 30282 7828 30288 7880
rect 30340 7828 30346 7880
rect 30300 7800 30328 7828
rect 27948 7772 30328 7800
rect 27948 7760 27954 7772
rect 25777 7735 25835 7741
rect 25777 7701 25789 7735
rect 25823 7732 25835 7735
rect 26326 7732 26332 7744
rect 25823 7704 26332 7732
rect 25823 7701 25835 7704
rect 25777 7695 25835 7701
rect 26326 7692 26332 7704
rect 26384 7692 26390 7744
rect 28261 7735 28319 7741
rect 28261 7701 28273 7735
rect 28307 7732 28319 7735
rect 28442 7732 28448 7744
rect 28307 7704 28448 7732
rect 28307 7701 28319 7704
rect 28261 7695 28319 7701
rect 28442 7692 28448 7704
rect 28500 7692 28506 7744
rect 1104 7642 38824 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 35594 7642
rect 35646 7590 35658 7642
rect 35710 7590 35722 7642
rect 35774 7590 35786 7642
rect 35838 7590 35850 7642
rect 35902 7590 38824 7642
rect 1104 7568 38824 7590
rect 22922 7488 22928 7540
rect 22980 7528 22986 7540
rect 24029 7531 24087 7537
rect 24029 7528 24041 7531
rect 22980 7500 24041 7528
rect 22980 7488 22986 7500
rect 24029 7497 24041 7500
rect 24075 7497 24087 7531
rect 24029 7491 24087 7497
rect 25866 7488 25872 7540
rect 25924 7528 25930 7540
rect 26973 7531 27031 7537
rect 26973 7528 26985 7531
rect 25924 7500 26985 7528
rect 25924 7488 25930 7500
rect 26973 7497 26985 7500
rect 27019 7497 27031 7531
rect 26973 7491 27031 7497
rect 28353 7531 28411 7537
rect 28353 7497 28365 7531
rect 28399 7528 28411 7531
rect 30190 7528 30196 7540
rect 28399 7500 30196 7528
rect 28399 7497 28411 7500
rect 28353 7491 28411 7497
rect 30190 7488 30196 7500
rect 30248 7488 30254 7540
rect 30282 7488 30288 7540
rect 30340 7488 30346 7540
rect 21269 7463 21327 7469
rect 21269 7460 21281 7463
rect 20732 7432 21281 7460
rect 20732 7401 20760 7432
rect 21269 7429 21281 7432
rect 21315 7429 21327 7463
rect 24486 7460 24492 7472
rect 21269 7423 21327 7429
rect 21468 7432 24492 7460
rect 21468 7401 21496 7432
rect 20717 7395 20775 7401
rect 20717 7361 20729 7395
rect 20763 7361 20775 7395
rect 20717 7355 20775 7361
rect 20993 7395 21051 7401
rect 20993 7361 21005 7395
rect 21039 7392 21051 7395
rect 21453 7395 21511 7401
rect 21453 7392 21465 7395
rect 21039 7364 21465 7392
rect 21039 7361 21051 7364
rect 20993 7355 21051 7361
rect 21453 7361 21465 7364
rect 21499 7361 21511 7395
rect 22005 7395 22063 7401
rect 22005 7392 22017 7395
rect 21453 7355 21511 7361
rect 21560 7364 22017 7392
rect 20809 7327 20867 7333
rect 20809 7293 20821 7327
rect 20855 7293 20867 7327
rect 20809 7287 20867 7293
rect 21177 7327 21235 7333
rect 21177 7293 21189 7327
rect 21223 7324 21235 7327
rect 21560 7324 21588 7364
rect 22005 7361 22017 7364
rect 22051 7361 22063 7395
rect 22005 7355 22063 7361
rect 23569 7395 23627 7401
rect 23569 7361 23581 7395
rect 23615 7361 23627 7395
rect 23569 7355 23627 7361
rect 21223 7296 21588 7324
rect 21637 7327 21695 7333
rect 21223 7293 21235 7296
rect 21177 7287 21235 7293
rect 21637 7293 21649 7327
rect 21683 7324 21695 7327
rect 22097 7327 22155 7333
rect 22097 7324 22109 7327
rect 21683 7296 22109 7324
rect 21683 7293 21695 7296
rect 21637 7287 21695 7293
rect 22097 7293 22109 7296
rect 22143 7293 22155 7327
rect 22097 7287 22155 7293
rect 20824 7256 20852 7287
rect 22738 7284 22744 7336
rect 22796 7324 22802 7336
rect 22796 7296 22968 7324
rect 22796 7284 22802 7296
rect 22833 7259 22891 7265
rect 22833 7256 22845 7259
rect 20824 7228 22845 7256
rect 22833 7225 22845 7228
rect 22879 7225 22891 7259
rect 22940 7256 22968 7296
rect 23014 7284 23020 7336
rect 23072 7324 23078 7336
rect 23477 7327 23535 7333
rect 23477 7324 23489 7327
rect 23072 7296 23489 7324
rect 23072 7284 23078 7296
rect 23477 7293 23489 7296
rect 23523 7324 23535 7327
rect 23584 7324 23612 7355
rect 23842 7352 23848 7404
rect 23900 7352 23906 7404
rect 24320 7401 24348 7432
rect 24486 7420 24492 7432
rect 24544 7420 24550 7472
rect 27890 7460 27896 7472
rect 27264 7432 27896 7460
rect 24305 7395 24363 7401
rect 24305 7361 24317 7395
rect 24351 7361 24363 7395
rect 24305 7355 24363 7361
rect 24394 7352 24400 7404
rect 24452 7352 24458 7404
rect 24765 7395 24823 7401
rect 24765 7361 24777 7395
rect 24811 7392 24823 7395
rect 24854 7392 24860 7404
rect 24811 7364 24860 7392
rect 24811 7361 24823 7364
rect 24765 7355 24823 7361
rect 24854 7352 24860 7364
rect 24912 7352 24918 7404
rect 26510 7352 26516 7404
rect 26568 7352 26574 7404
rect 26602 7352 26608 7404
rect 26660 7352 26666 7404
rect 26789 7395 26847 7401
rect 26789 7361 26801 7395
rect 26835 7392 26847 7395
rect 26970 7392 26976 7404
rect 26835 7364 26976 7392
rect 26835 7361 26847 7364
rect 26789 7355 26847 7361
rect 26970 7352 26976 7364
rect 27028 7352 27034 7404
rect 27264 7401 27292 7432
rect 27890 7420 27896 7432
rect 27948 7420 27954 7472
rect 28902 7460 28908 7472
rect 28552 7432 28908 7460
rect 27249 7395 27307 7401
rect 27249 7361 27261 7395
rect 27295 7361 27307 7395
rect 27249 7355 27307 7361
rect 27433 7395 27491 7401
rect 27433 7361 27445 7395
rect 27479 7390 27491 7395
rect 27614 7392 27620 7404
rect 27540 7390 27620 7392
rect 27479 7364 27620 7390
rect 27479 7362 27568 7364
rect 27479 7361 27491 7362
rect 27433 7355 27491 7361
rect 27614 7352 27620 7364
rect 27672 7392 27678 7404
rect 27672 7364 28120 7392
rect 27672 7352 27678 7364
rect 23523 7296 23612 7324
rect 23523 7293 23535 7296
rect 23477 7287 23535 7293
rect 23658 7284 23664 7336
rect 23716 7284 23722 7336
rect 27154 7284 27160 7336
rect 27212 7284 27218 7336
rect 27338 7284 27344 7336
rect 27396 7284 27402 7336
rect 27798 7284 27804 7336
rect 27856 7284 27862 7336
rect 27890 7284 27896 7336
rect 27948 7284 27954 7336
rect 28092 7333 28120 7364
rect 28258 7352 28264 7404
rect 28316 7352 28322 7404
rect 28442 7352 28448 7404
rect 28500 7352 28506 7404
rect 28552 7401 28580 7432
rect 28902 7420 28908 7432
rect 28960 7460 28966 7472
rect 29086 7460 29092 7472
rect 28960 7432 29092 7460
rect 28960 7420 28966 7432
rect 29086 7420 29092 7432
rect 29144 7420 29150 7472
rect 29270 7420 29276 7472
rect 29328 7420 29334 7472
rect 28537 7395 28595 7401
rect 28537 7361 28549 7395
rect 28583 7361 28595 7395
rect 28537 7355 28595 7361
rect 29822 7352 29828 7404
rect 29880 7352 29886 7404
rect 27985 7327 28043 7333
rect 27985 7293 27997 7327
rect 28031 7293 28043 7327
rect 27985 7287 28043 7293
rect 28077 7327 28135 7333
rect 28077 7293 28089 7327
rect 28123 7293 28135 7327
rect 28077 7287 28135 7293
rect 22940 7228 23612 7256
rect 22833 7219 22891 7225
rect 20530 7148 20536 7200
rect 20588 7148 20594 7200
rect 21818 7148 21824 7200
rect 21876 7148 21882 7200
rect 23584 7197 23612 7228
rect 27522 7216 27528 7268
rect 27580 7256 27586 7268
rect 27617 7259 27675 7265
rect 27617 7256 27629 7259
rect 27580 7228 27629 7256
rect 27580 7216 27586 7228
rect 27617 7225 27629 7228
rect 27663 7225 27675 7259
rect 27617 7219 27675 7225
rect 28000 7256 28028 7287
rect 28350 7256 28356 7268
rect 28000 7228 28356 7256
rect 23569 7191 23627 7197
rect 23569 7157 23581 7191
rect 23615 7157 23627 7191
rect 23569 7151 23627 7157
rect 24118 7148 24124 7200
rect 24176 7148 24182 7200
rect 24302 7148 24308 7200
rect 24360 7188 24366 7200
rect 24581 7191 24639 7197
rect 24581 7188 24593 7191
rect 24360 7160 24593 7188
rect 24360 7148 24366 7160
rect 24581 7157 24593 7160
rect 24627 7157 24639 7191
rect 24581 7151 24639 7157
rect 26694 7148 26700 7200
rect 26752 7148 26758 7200
rect 27338 7148 27344 7200
rect 27396 7188 27402 7200
rect 28000 7188 28028 7228
rect 28350 7216 28356 7228
rect 28408 7216 28414 7268
rect 27396 7160 28028 7188
rect 28460 7188 28488 7352
rect 28813 7327 28871 7333
rect 28813 7293 28825 7327
rect 28859 7324 28871 7327
rect 29840 7324 29868 7352
rect 28859 7296 29868 7324
rect 28859 7293 28871 7296
rect 28813 7287 28871 7293
rect 28902 7188 28908 7200
rect 28460 7160 28908 7188
rect 27396 7148 27402 7160
rect 28902 7148 28908 7160
rect 28960 7148 28966 7200
rect 1104 7098 38824 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38824 7098
rect 1104 7024 38824 7046
rect 20428 6987 20486 6993
rect 20428 6953 20440 6987
rect 20474 6984 20486 6987
rect 20530 6984 20536 6996
rect 20474 6956 20536 6984
rect 20474 6953 20486 6956
rect 20428 6947 20486 6953
rect 20530 6944 20536 6956
rect 20588 6944 20594 6996
rect 24854 6944 24860 6996
rect 24912 6944 24918 6996
rect 26694 6984 26700 6996
rect 25884 6956 26700 6984
rect 23492 6888 23888 6916
rect 23492 6860 23520 6888
rect 23860 6860 23888 6888
rect 20165 6851 20223 6857
rect 20165 6817 20177 6851
rect 20211 6848 20223 6851
rect 20806 6848 20812 6860
rect 20211 6820 20812 6848
rect 20211 6817 20223 6820
rect 20165 6811 20223 6817
rect 20806 6808 20812 6820
rect 20864 6808 20870 6860
rect 21913 6851 21971 6857
rect 21913 6817 21925 6851
rect 21959 6848 21971 6851
rect 22738 6848 22744 6860
rect 21959 6820 22744 6848
rect 21959 6817 21971 6820
rect 21913 6811 21971 6817
rect 22738 6808 22744 6820
rect 22796 6808 22802 6860
rect 23474 6848 23480 6860
rect 22873 6820 23480 6848
rect 22186 6780 22192 6792
rect 21574 6752 22192 6780
rect 22186 6740 22192 6752
rect 22244 6780 22250 6792
rect 22465 6783 22523 6789
rect 22465 6780 22477 6783
rect 22244 6752 22477 6780
rect 22244 6740 22250 6752
rect 22465 6749 22477 6752
rect 22511 6780 22523 6783
rect 22554 6780 22560 6792
rect 22511 6752 22560 6780
rect 22511 6749 22523 6752
rect 22465 6743 22523 6749
rect 22554 6740 22560 6752
rect 22612 6740 22618 6792
rect 22649 6783 22707 6789
rect 22649 6749 22661 6783
rect 22695 6780 22707 6783
rect 22873 6780 22901 6820
rect 23474 6808 23480 6820
rect 23532 6808 23538 6860
rect 23658 6808 23664 6860
rect 23716 6808 23722 6860
rect 23842 6808 23848 6860
rect 23900 6808 23906 6860
rect 24213 6851 24271 6857
rect 24213 6817 24225 6851
rect 24259 6848 24271 6851
rect 24765 6851 24823 6857
rect 24765 6848 24777 6851
rect 24259 6820 24777 6848
rect 24259 6817 24271 6820
rect 24213 6811 24271 6817
rect 24765 6817 24777 6820
rect 24811 6817 24823 6851
rect 24765 6811 24823 6817
rect 25409 6851 25467 6857
rect 25409 6817 25421 6851
rect 25455 6817 25467 6851
rect 25409 6811 25467 6817
rect 22695 6752 22901 6780
rect 23293 6783 23351 6789
rect 22695 6749 22707 6752
rect 22649 6743 22707 6749
rect 23293 6749 23305 6783
rect 23339 6780 23351 6783
rect 24118 6780 24124 6792
rect 23339 6752 24124 6780
rect 23339 6749 23351 6752
rect 23293 6743 23351 6749
rect 24118 6740 24124 6752
rect 24176 6740 24182 6792
rect 24394 6740 24400 6792
rect 24452 6740 24458 6792
rect 24486 6740 24492 6792
rect 24544 6780 24550 6792
rect 24581 6783 24639 6789
rect 24581 6780 24593 6783
rect 24544 6752 24593 6780
rect 24544 6740 24550 6752
rect 24581 6749 24593 6752
rect 24627 6780 24639 6783
rect 25317 6783 25375 6789
rect 25317 6780 25329 6783
rect 24627 6752 25329 6780
rect 24627 6749 24639 6752
rect 24581 6743 24639 6749
rect 25317 6749 25329 6752
rect 25363 6749 25375 6783
rect 25424 6780 25452 6811
rect 25498 6780 25504 6792
rect 25424 6752 25504 6780
rect 25317 6743 25375 6749
rect 25498 6740 25504 6752
rect 25556 6740 25562 6792
rect 25884 6789 25912 6956
rect 26694 6944 26700 6956
rect 26752 6944 26758 6996
rect 26973 6987 27031 6993
rect 26973 6953 26985 6987
rect 27019 6984 27031 6987
rect 27798 6984 27804 6996
rect 27019 6956 27804 6984
rect 27019 6953 27031 6956
rect 26973 6947 27031 6953
rect 27798 6944 27804 6956
rect 27856 6984 27862 6996
rect 27893 6987 27951 6993
rect 27893 6984 27905 6987
rect 27856 6956 27905 6984
rect 27856 6944 27862 6956
rect 27893 6953 27905 6956
rect 27939 6953 27951 6987
rect 27893 6947 27951 6953
rect 28626 6944 28632 6996
rect 28684 6944 28690 6996
rect 28810 6944 28816 6996
rect 28868 6984 28874 6996
rect 29549 6987 29607 6993
rect 29549 6984 29561 6987
rect 28868 6956 29561 6984
rect 28868 6944 28874 6956
rect 29549 6953 29561 6956
rect 29595 6984 29607 6987
rect 29730 6984 29736 6996
rect 29595 6956 29736 6984
rect 29595 6953 29607 6956
rect 29549 6947 29607 6953
rect 29730 6944 29736 6956
rect 29788 6944 29794 6996
rect 29825 6987 29883 6993
rect 29825 6953 29837 6987
rect 29871 6984 29883 6987
rect 30006 6984 30012 6996
rect 29871 6956 30012 6984
rect 29871 6953 29883 6956
rect 29825 6947 29883 6953
rect 30006 6944 30012 6956
rect 30064 6944 30070 6996
rect 26326 6876 26332 6928
rect 26384 6876 26390 6928
rect 27154 6876 27160 6928
rect 27212 6916 27218 6928
rect 28997 6919 29055 6925
rect 28997 6916 29009 6919
rect 27212 6888 27752 6916
rect 27212 6876 27218 6888
rect 26344 6848 26372 6876
rect 27724 6848 27752 6888
rect 28736 6888 29009 6916
rect 28736 6848 28764 6888
rect 28997 6885 29009 6888
rect 29043 6885 29055 6919
rect 28997 6879 29055 6885
rect 26206 6820 26372 6848
rect 26620 6820 27292 6848
rect 27724 6820 28764 6848
rect 25869 6783 25927 6789
rect 25869 6749 25881 6783
rect 25915 6749 25927 6783
rect 25869 6743 25927 6749
rect 26050 6740 26056 6792
rect 26108 6740 26114 6792
rect 26206 6789 26234 6820
rect 26620 6792 26648 6820
rect 26191 6783 26249 6789
rect 26191 6749 26203 6783
rect 26237 6749 26249 6783
rect 26191 6743 26249 6749
rect 26326 6740 26332 6792
rect 26384 6740 26390 6792
rect 26421 6783 26479 6789
rect 26421 6749 26433 6783
rect 26467 6749 26479 6783
rect 26421 6743 26479 6749
rect 22094 6672 22100 6724
rect 22152 6712 22158 6724
rect 23106 6712 23112 6724
rect 22152 6684 23112 6712
rect 22152 6672 22158 6684
rect 23106 6672 23112 6684
rect 23164 6672 23170 6724
rect 23201 6715 23259 6721
rect 23201 6681 23213 6715
rect 23247 6712 23259 6715
rect 24412 6712 24440 6740
rect 23247 6684 24440 6712
rect 25225 6715 25283 6721
rect 23247 6681 23259 6684
rect 23201 6675 23259 6681
rect 25225 6681 25237 6715
rect 25271 6712 25283 6715
rect 25961 6715 26019 6721
rect 25271 6684 25912 6712
rect 25271 6681 25283 6684
rect 25225 6675 25283 6681
rect 20714 6604 20720 6656
rect 20772 6644 20778 6656
rect 21818 6644 21824 6656
rect 20772 6616 21824 6644
rect 20772 6604 20778 6616
rect 21818 6604 21824 6616
rect 21876 6604 21882 6656
rect 23477 6647 23535 6653
rect 23477 6613 23489 6647
rect 23523 6644 23535 6647
rect 23658 6644 23664 6656
rect 23523 6616 23664 6644
rect 23523 6613 23535 6616
rect 23477 6607 23535 6613
rect 23658 6604 23664 6616
rect 23716 6604 23722 6656
rect 24394 6604 24400 6656
rect 24452 6604 24458 6656
rect 25682 6604 25688 6656
rect 25740 6604 25746 6656
rect 25884 6644 25912 6684
rect 25961 6681 25973 6715
rect 26007 6712 26019 6715
rect 26436 6712 26464 6743
rect 26602 6740 26608 6792
rect 26660 6740 26666 6792
rect 26881 6783 26939 6789
rect 26881 6749 26893 6783
rect 26927 6780 26939 6783
rect 26970 6780 26976 6792
rect 26927 6752 26976 6780
rect 26927 6749 26939 6752
rect 26881 6743 26939 6749
rect 26970 6740 26976 6752
rect 27028 6740 27034 6792
rect 27264 6789 27292 6820
rect 28902 6808 28908 6860
rect 28960 6848 28966 6860
rect 28960 6820 29868 6848
rect 28960 6808 28966 6820
rect 27249 6783 27307 6789
rect 27249 6749 27261 6783
rect 27295 6749 27307 6783
rect 27249 6743 27307 6749
rect 27341 6783 27399 6789
rect 27341 6749 27353 6783
rect 27387 6780 27399 6783
rect 27430 6780 27436 6792
rect 27387 6752 27436 6780
rect 27387 6749 27399 6752
rect 27341 6743 27399 6749
rect 26007 6684 26464 6712
rect 26007 6681 26019 6684
rect 25961 6675 26019 6681
rect 26510 6672 26516 6724
rect 26568 6712 26574 6724
rect 26789 6715 26847 6721
rect 26789 6712 26801 6715
rect 26568 6684 26801 6712
rect 26568 6672 26574 6684
rect 26789 6681 26801 6684
rect 26835 6712 26847 6715
rect 27356 6712 27384 6743
rect 27430 6740 27436 6752
rect 27488 6740 27494 6792
rect 27614 6740 27620 6792
rect 27672 6740 27678 6792
rect 27706 6740 27712 6792
rect 27764 6780 27770 6792
rect 27801 6783 27859 6789
rect 27801 6780 27813 6783
rect 27764 6752 27813 6780
rect 27764 6740 27770 6752
rect 27801 6749 27813 6752
rect 27847 6749 27859 6783
rect 28320 6783 28378 6789
rect 28320 6780 28332 6783
rect 27801 6743 27859 6749
rect 28000 6752 28332 6780
rect 26835 6684 27384 6712
rect 27525 6715 27583 6721
rect 26835 6681 26847 6684
rect 26789 6675 26847 6681
rect 27525 6681 27537 6715
rect 27571 6712 27583 6715
rect 27632 6712 27660 6740
rect 28000 6712 28028 6752
rect 28320 6749 28332 6752
rect 28366 6749 28378 6783
rect 28320 6743 28378 6749
rect 28442 6740 28448 6792
rect 28500 6780 28506 6792
rect 28552 6789 28764 6790
rect 29840 6789 29868 6820
rect 28552 6783 28779 6789
rect 28552 6780 28733 6783
rect 28500 6762 28733 6780
rect 28500 6752 28580 6762
rect 28500 6740 28506 6752
rect 28721 6749 28733 6762
rect 28767 6749 28779 6783
rect 28721 6743 28779 6749
rect 28813 6783 28871 6789
rect 28813 6749 28825 6783
rect 28859 6749 28871 6783
rect 28813 6743 28871 6749
rect 29825 6783 29883 6789
rect 29825 6749 29837 6783
rect 29871 6749 29883 6783
rect 29825 6743 29883 6749
rect 30009 6783 30067 6789
rect 30009 6749 30021 6783
rect 30055 6749 30067 6783
rect 30009 6743 30067 6749
rect 28537 6715 28595 6721
rect 28537 6712 28549 6715
rect 27571 6684 28028 6712
rect 28092 6684 28549 6712
rect 27571 6681 27583 6684
rect 27525 6675 27583 6681
rect 26050 6644 26056 6656
rect 25884 6616 26056 6644
rect 26050 6604 26056 6616
rect 26108 6604 26114 6656
rect 26970 6604 26976 6656
rect 27028 6644 27034 6656
rect 27157 6647 27215 6653
rect 27157 6644 27169 6647
rect 27028 6616 27169 6644
rect 27028 6604 27034 6616
rect 27157 6613 27169 6616
rect 27203 6644 27215 6647
rect 27430 6644 27436 6656
rect 27203 6616 27436 6644
rect 27203 6613 27215 6616
rect 27157 6607 27215 6613
rect 27430 6604 27436 6616
rect 27488 6644 27494 6656
rect 28092 6644 28120 6684
rect 28537 6681 28549 6684
rect 28583 6681 28595 6715
rect 28537 6675 28595 6681
rect 28828 6656 28856 6743
rect 28902 6672 28908 6724
rect 28960 6712 28966 6724
rect 30024 6712 30052 6743
rect 28960 6684 30052 6712
rect 28960 6672 28966 6684
rect 27488 6616 28120 6644
rect 28261 6647 28319 6653
rect 27488 6604 27494 6616
rect 28261 6613 28273 6647
rect 28307 6644 28319 6647
rect 28350 6644 28356 6656
rect 28307 6616 28356 6644
rect 28307 6613 28319 6616
rect 28261 6607 28319 6613
rect 28350 6604 28356 6616
rect 28408 6604 28414 6656
rect 28442 6604 28448 6656
rect 28500 6604 28506 6656
rect 28810 6604 28816 6656
rect 28868 6604 28874 6656
rect 1104 6554 38824 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 35594 6554
rect 35646 6502 35658 6554
rect 35710 6502 35722 6554
rect 35774 6502 35786 6554
rect 35838 6502 35850 6554
rect 35902 6502 38824 6554
rect 1104 6480 38824 6502
rect 20806 6440 20812 6452
rect 19904 6412 20812 6440
rect 19904 6313 19932 6412
rect 20806 6400 20812 6412
rect 20864 6400 20870 6452
rect 21637 6443 21695 6449
rect 21637 6409 21649 6443
rect 21683 6440 21695 6443
rect 23014 6440 23020 6452
rect 21683 6412 23020 6440
rect 21683 6409 21695 6412
rect 21637 6403 21695 6409
rect 23014 6400 23020 6412
rect 23072 6400 23078 6452
rect 23106 6400 23112 6452
rect 23164 6440 23170 6452
rect 23164 6412 23520 6440
rect 23164 6400 23170 6412
rect 22186 6372 22192 6384
rect 21390 6344 22192 6372
rect 22186 6332 22192 6344
rect 22244 6372 22250 6384
rect 22646 6372 22652 6384
rect 22244 6344 22652 6372
rect 22244 6332 22250 6344
rect 22646 6332 22652 6344
rect 22704 6332 22710 6384
rect 23492 6372 23520 6412
rect 23566 6400 23572 6452
rect 23624 6440 23630 6452
rect 23661 6443 23719 6449
rect 23661 6440 23673 6443
rect 23624 6412 23673 6440
rect 23624 6400 23630 6412
rect 23661 6409 23673 6412
rect 23707 6409 23719 6443
rect 23661 6403 23719 6409
rect 23768 6412 25360 6440
rect 23768 6372 23796 6412
rect 25332 6384 25360 6412
rect 25498 6400 25504 6452
rect 25556 6400 25562 6452
rect 25774 6400 25780 6452
rect 25832 6440 25838 6452
rect 25869 6443 25927 6449
rect 25869 6440 25881 6443
rect 25832 6412 25881 6440
rect 25832 6400 25838 6412
rect 25869 6409 25881 6412
rect 25915 6409 25927 6443
rect 25869 6403 25927 6409
rect 26326 6400 26332 6452
rect 26384 6440 26390 6452
rect 26973 6443 27031 6449
rect 26973 6440 26985 6443
rect 26384 6412 26985 6440
rect 26384 6400 26390 6412
rect 26973 6409 26985 6412
rect 27019 6409 27031 6443
rect 26973 6403 27031 6409
rect 27614 6400 27620 6452
rect 27672 6440 27678 6452
rect 27709 6443 27767 6449
rect 27709 6440 27721 6443
rect 27672 6412 27721 6440
rect 27672 6400 27678 6412
rect 27709 6409 27721 6412
rect 27755 6440 27767 6443
rect 28810 6440 28816 6452
rect 27755 6412 28816 6440
rect 27755 6409 27767 6412
rect 27709 6403 27767 6409
rect 28810 6400 28816 6412
rect 28868 6400 28874 6452
rect 29086 6400 29092 6452
rect 29144 6400 29150 6452
rect 23492 6344 23796 6372
rect 24029 6375 24087 6381
rect 24029 6341 24041 6375
rect 24075 6372 24087 6375
rect 24302 6372 24308 6384
rect 24075 6344 24308 6372
rect 24075 6341 24087 6344
rect 24029 6335 24087 6341
rect 24302 6332 24308 6344
rect 24360 6332 24366 6384
rect 25314 6332 25320 6384
rect 25372 6332 25378 6384
rect 25516 6372 25544 6400
rect 25516 6344 26832 6372
rect 19889 6307 19947 6313
rect 19889 6273 19901 6307
rect 19935 6273 19947 6307
rect 25332 6304 25360 6332
rect 25777 6307 25835 6313
rect 25777 6304 25789 6307
rect 19889 6267 19947 6273
rect 20165 6239 20223 6245
rect 20165 6205 20177 6239
rect 20211 6236 20223 6239
rect 20714 6236 20720 6248
rect 20211 6208 20720 6236
rect 20211 6205 20223 6208
rect 20165 6199 20223 6205
rect 20714 6196 20720 6208
rect 20772 6196 20778 6248
rect 20806 6196 20812 6248
rect 20864 6236 20870 6248
rect 21913 6239 21971 6245
rect 21913 6236 21925 6239
rect 20864 6208 21925 6236
rect 20864 6196 20870 6208
rect 21913 6205 21925 6208
rect 21959 6205 21971 6239
rect 21913 6199 21971 6205
rect 21928 6100 21956 6199
rect 22186 6196 22192 6248
rect 22244 6196 22250 6248
rect 23753 6239 23811 6245
rect 23753 6236 23765 6239
rect 23584 6208 23765 6236
rect 23584 6112 23612 6208
rect 23753 6205 23765 6208
rect 23799 6205 23811 6239
rect 25148 6236 25176 6290
rect 25332 6276 25789 6304
rect 25777 6273 25789 6276
rect 25823 6273 25835 6307
rect 25777 6267 25835 6273
rect 26602 6264 26608 6316
rect 26660 6264 26666 6316
rect 26804 6313 26832 6344
rect 27890 6332 27896 6384
rect 27948 6372 27954 6384
rect 29104 6372 29132 6400
rect 27948 6344 28014 6372
rect 29104 6344 29500 6372
rect 27948 6332 27954 6344
rect 26789 6307 26847 6313
rect 26789 6273 26801 6307
rect 26835 6304 26847 6307
rect 27430 6304 27436 6316
rect 26835 6276 27436 6304
rect 26835 6273 26847 6276
rect 26789 6267 26847 6273
rect 27430 6264 27436 6276
rect 27488 6264 27494 6316
rect 29472 6313 29500 6344
rect 29457 6307 29515 6313
rect 29457 6273 29469 6307
rect 29503 6273 29515 6307
rect 29457 6267 29515 6273
rect 26513 6239 26571 6245
rect 25148 6208 25820 6236
rect 23753 6199 23811 6205
rect 25792 6180 25820 6208
rect 26513 6205 26525 6239
rect 26559 6205 26571 6239
rect 26620 6236 26648 6264
rect 27525 6239 27583 6245
rect 27525 6236 27537 6239
rect 26620 6208 27537 6236
rect 26513 6199 26571 6205
rect 27525 6205 27537 6208
rect 27571 6236 27583 6239
rect 28534 6236 28540 6248
rect 27571 6208 28540 6236
rect 27571 6205 27583 6208
rect 27525 6199 27583 6205
rect 25774 6128 25780 6180
rect 25832 6128 25838 6180
rect 26528 6168 26556 6199
rect 28534 6196 28540 6208
rect 28592 6196 28598 6248
rect 29086 6196 29092 6248
rect 29144 6236 29150 6248
rect 29181 6239 29239 6245
rect 29181 6236 29193 6239
rect 29144 6208 29193 6236
rect 29144 6196 29150 6208
rect 29181 6205 29193 6208
rect 29227 6205 29239 6239
rect 29181 6199 29239 6205
rect 27154 6168 27160 6180
rect 26528 6140 27160 6168
rect 27154 6128 27160 6140
rect 27212 6168 27218 6180
rect 27706 6168 27712 6180
rect 27212 6140 27712 6168
rect 27212 6128 27218 6140
rect 27706 6128 27712 6140
rect 27764 6128 27770 6180
rect 23566 6100 23572 6112
rect 21928 6072 23572 6100
rect 23566 6060 23572 6072
rect 23624 6060 23630 6112
rect 26234 6060 26240 6112
rect 26292 6060 26298 6112
rect 26510 6060 26516 6112
rect 26568 6060 26574 6112
rect 1104 6010 38824 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38824 6010
rect 1104 5936 38824 5958
rect 22189 5899 22247 5905
rect 22189 5865 22201 5899
rect 22235 5896 22247 5899
rect 23474 5896 23480 5908
rect 22235 5868 23480 5896
rect 22235 5865 22247 5868
rect 22189 5859 22247 5865
rect 23474 5856 23480 5868
rect 23532 5856 23538 5908
rect 23566 5856 23572 5908
rect 23624 5896 23630 5908
rect 23624 5868 23980 5896
rect 23624 5856 23630 5868
rect 23658 5720 23664 5772
rect 23716 5720 23722 5772
rect 23952 5769 23980 5868
rect 25682 5856 25688 5908
rect 25740 5856 25746 5908
rect 26145 5899 26203 5905
rect 26145 5865 26157 5899
rect 26191 5896 26203 5899
rect 26602 5896 26608 5908
rect 26191 5868 26608 5896
rect 26191 5865 26203 5868
rect 26145 5859 26203 5865
rect 26602 5856 26608 5868
rect 26660 5856 26666 5908
rect 27982 5856 27988 5908
rect 28040 5856 28046 5908
rect 28442 5856 28448 5908
rect 28500 5856 28506 5908
rect 28905 5899 28963 5905
rect 28905 5865 28917 5899
rect 28951 5896 28963 5899
rect 29086 5896 29092 5908
rect 28951 5868 29092 5896
rect 28951 5865 28963 5868
rect 28905 5859 28963 5865
rect 29086 5856 29092 5868
rect 29144 5856 29150 5908
rect 23937 5763 23995 5769
rect 23937 5729 23949 5763
rect 23983 5760 23995 5763
rect 24397 5763 24455 5769
rect 24397 5760 24409 5763
rect 23983 5732 24409 5760
rect 23983 5729 23995 5732
rect 23937 5723 23995 5729
rect 24397 5729 24409 5732
rect 24443 5729 24455 5763
rect 24397 5723 24455 5729
rect 24673 5763 24731 5769
rect 24673 5729 24685 5763
rect 24719 5760 24731 5763
rect 25700 5760 25728 5856
rect 24719 5732 25728 5760
rect 26237 5763 26295 5769
rect 24719 5729 24731 5732
rect 24673 5723 24731 5729
rect 26237 5729 26249 5763
rect 26283 5760 26295 5763
rect 27062 5760 27068 5772
rect 26283 5732 27068 5760
rect 26283 5729 26295 5732
rect 26237 5723 26295 5729
rect 27062 5720 27068 5732
rect 27120 5720 27126 5772
rect 28460 5760 28488 5856
rect 28460 5732 28948 5760
rect 22646 5692 22652 5704
rect 22586 5664 22652 5692
rect 22646 5652 22652 5664
rect 22704 5652 22710 5704
rect 25774 5652 25780 5704
rect 25832 5652 25838 5704
rect 27890 5692 27896 5704
rect 27646 5664 27896 5692
rect 27890 5652 27896 5664
rect 27948 5652 27954 5704
rect 28810 5652 28816 5704
rect 28868 5652 28874 5704
rect 28920 5701 28948 5732
rect 28905 5695 28963 5701
rect 28905 5661 28917 5695
rect 28951 5661 28963 5695
rect 28905 5655 28963 5661
rect 29181 5695 29239 5701
rect 29181 5661 29193 5695
rect 29227 5661 29239 5695
rect 29181 5655 29239 5661
rect 26510 5584 26516 5636
rect 26568 5584 26574 5636
rect 29196 5624 29224 5655
rect 27816 5596 29224 5624
rect 26694 5516 26700 5568
rect 26752 5556 26758 5568
rect 27816 5556 27844 5596
rect 26752 5528 27844 5556
rect 26752 5516 26758 5528
rect 28166 5516 28172 5568
rect 28224 5516 28230 5568
rect 29086 5516 29092 5568
rect 29144 5516 29150 5568
rect 1104 5466 38824 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 35594 5466
rect 35646 5414 35658 5466
rect 35710 5414 35722 5466
rect 35774 5414 35786 5466
rect 35838 5414 35850 5466
rect 35902 5414 38824 5466
rect 1104 5392 38824 5414
rect 22186 5312 22192 5364
rect 22244 5352 22250 5364
rect 22465 5355 22523 5361
rect 22465 5352 22477 5355
rect 22244 5324 22477 5352
rect 22244 5312 22250 5324
rect 22465 5321 22477 5324
rect 22511 5321 22523 5355
rect 22465 5315 22523 5321
rect 24394 5312 24400 5364
rect 24452 5312 24458 5364
rect 25961 5355 26019 5361
rect 25961 5321 25973 5355
rect 26007 5352 26019 5355
rect 26234 5352 26240 5364
rect 26007 5324 26240 5352
rect 26007 5321 26019 5324
rect 25961 5315 26019 5321
rect 26234 5312 26240 5324
rect 26292 5312 26298 5364
rect 26510 5312 26516 5364
rect 26568 5352 26574 5364
rect 26605 5355 26663 5361
rect 26605 5352 26617 5355
rect 26568 5324 26617 5352
rect 26568 5312 26574 5324
rect 26605 5321 26617 5324
rect 26651 5321 26663 5355
rect 26605 5315 26663 5321
rect 28166 5312 28172 5364
rect 28224 5312 28230 5364
rect 28537 5355 28595 5361
rect 28537 5321 28549 5355
rect 28583 5352 28595 5355
rect 29086 5352 29092 5364
rect 28583 5324 29092 5352
rect 28583 5321 28595 5324
rect 28537 5315 28595 5321
rect 29086 5312 29092 5324
rect 29144 5312 29150 5364
rect 22649 5219 22707 5225
rect 22649 5185 22661 5219
rect 22695 5216 22707 5219
rect 24412 5216 24440 5312
rect 22695 5188 24440 5216
rect 26329 5219 26387 5225
rect 22695 5185 22707 5188
rect 22649 5179 22707 5185
rect 26329 5185 26341 5219
rect 26375 5216 26387 5219
rect 27157 5219 27215 5225
rect 27157 5216 27169 5219
rect 26375 5188 27169 5216
rect 26375 5185 26387 5188
rect 26329 5179 26387 5185
rect 27157 5185 27169 5188
rect 27203 5185 27215 5219
rect 27157 5179 27215 5185
rect 27801 5219 27859 5225
rect 27801 5185 27813 5219
rect 27847 5216 27859 5219
rect 27982 5216 27988 5228
rect 27847 5188 27988 5216
rect 27847 5185 27859 5188
rect 27801 5179 27859 5185
rect 27982 5176 27988 5188
rect 28040 5176 28046 5228
rect 28184 5216 28212 5312
rect 28445 5219 28503 5225
rect 28445 5216 28457 5219
rect 28184 5188 28457 5216
rect 28445 5185 28457 5188
rect 28491 5185 28503 5219
rect 28445 5179 28503 5185
rect 26418 5108 26424 5160
rect 26476 5108 26482 5160
rect 1104 4922 38824 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38824 4922
rect 1104 4848 38824 4870
rect 26418 4768 26424 4820
rect 26476 4808 26482 4820
rect 27249 4811 27307 4817
rect 27249 4808 27261 4811
rect 26476 4780 27261 4808
rect 26476 4768 26482 4780
rect 27249 4777 27261 4780
rect 27295 4777 27307 4811
rect 27249 4771 27307 4777
rect 28350 4768 28356 4820
rect 28408 4768 28414 4820
rect 26973 4743 27031 4749
rect 26973 4709 26985 4743
rect 27019 4740 27031 4743
rect 28368 4740 28396 4768
rect 27019 4712 28396 4740
rect 27019 4709 27031 4712
rect 26973 4703 27031 4709
rect 27154 4564 27160 4616
rect 27212 4604 27218 4616
rect 27249 4607 27307 4613
rect 27249 4604 27261 4607
rect 27212 4576 27261 4604
rect 27212 4564 27218 4576
rect 27249 4573 27261 4576
rect 27295 4573 27307 4607
rect 27249 4567 27307 4573
rect 27430 4564 27436 4616
rect 27488 4564 27494 4616
rect 1104 4378 38824 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 35594 4378
rect 35646 4326 35658 4378
rect 35710 4326 35722 4378
rect 35774 4326 35786 4378
rect 35838 4326 35850 4378
rect 35902 4326 38824 4378
rect 1104 4304 38824 4326
rect 1104 3834 38824 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38824 3834
rect 1104 3760 38824 3782
rect 1104 3290 38824 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 35594 3290
rect 35646 3238 35658 3290
rect 35710 3238 35722 3290
rect 35774 3238 35786 3290
rect 35838 3238 35850 3290
rect 35902 3238 38824 3290
rect 1104 3216 38824 3238
rect 1104 2746 38824 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38824 2746
rect 1104 2672 38824 2694
rect 23937 2635 23995 2641
rect 23937 2601 23949 2635
rect 23983 2632 23995 2635
rect 24210 2632 24216 2644
rect 23983 2604 24216 2632
rect 23983 2601 23995 2604
rect 23937 2595 23995 2601
rect 24210 2592 24216 2604
rect 24268 2592 24274 2644
rect 23842 2388 23848 2440
rect 23900 2428 23906 2440
rect 24121 2431 24179 2437
rect 24121 2428 24133 2431
rect 23900 2400 24133 2428
rect 23900 2388 23906 2400
rect 24121 2397 24133 2400
rect 24167 2397 24179 2431
rect 24121 2391 24179 2397
rect 14 2320 20 2372
rect 72 2360 78 2372
rect 1489 2363 1547 2369
rect 1489 2360 1501 2363
rect 72 2332 1501 2360
rect 72 2320 78 2332
rect 1489 2329 1501 2332
rect 1535 2329 1547 2363
rect 1489 2323 1547 2329
rect 1673 2363 1731 2369
rect 1673 2329 1685 2363
rect 1719 2360 1731 2363
rect 1719 2332 6914 2360
rect 1719 2329 1731 2332
rect 1673 2323 1731 2329
rect 6886 2292 6914 2332
rect 11790 2320 11796 2372
rect 11848 2320 11854 2372
rect 11977 2363 12035 2369
rect 11977 2329 11989 2363
rect 12023 2360 12035 2363
rect 22094 2360 22100 2372
rect 12023 2332 22100 2360
rect 12023 2329 12035 2332
rect 11977 2323 12035 2329
rect 22094 2320 22100 2332
rect 22152 2320 22158 2372
rect 35529 2363 35587 2369
rect 35529 2360 35541 2363
rect 26206 2332 35541 2360
rect 18690 2292 18696 2304
rect 6886 2264 18696 2292
rect 18690 2252 18696 2264
rect 18748 2252 18754 2304
rect 22002 2252 22008 2304
rect 22060 2292 22066 2304
rect 26206 2292 26234 2332
rect 35529 2329 35541 2332
rect 35575 2329 35587 2363
rect 35529 2323 35587 2329
rect 35713 2363 35771 2369
rect 35713 2329 35725 2363
rect 35759 2329 35771 2363
rect 35713 2323 35771 2329
rect 22060 2264 26234 2292
rect 22060 2252 22066 2264
rect 35434 2252 35440 2304
rect 35492 2292 35498 2304
rect 35728 2292 35756 2323
rect 35492 2264 35756 2292
rect 35492 2252 35498 2264
rect 1104 2202 38824 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 35594 2202
rect 35646 2150 35658 2202
rect 35710 2150 35722 2202
rect 35774 2150 35786 2202
rect 35838 2150 35850 2202
rect 35902 2150 38824 2202
rect 1104 2128 38824 2150
<< via1 >>
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 940 37408 992 37460
rect 9680 37408 9732 37460
rect 21916 37272 21968 37324
rect 22284 37247 22336 37256
rect 22284 37213 22293 37247
rect 22293 37213 22327 37247
rect 22327 37213 22336 37247
rect 22284 37204 22336 37213
rect 33508 37204 33560 37256
rect 10140 37179 10192 37188
rect 10140 37145 10149 37179
rect 10149 37145 10183 37179
rect 10183 37145 10192 37179
rect 10140 37136 10192 37145
rect 26240 37136 26292 37188
rect 33692 37111 33744 37120
rect 33692 37077 33701 37111
rect 33701 37077 33735 37111
rect 33735 37077 33744 37111
rect 33692 37068 33744 37077
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 35594 36966 35646 37018
rect 35658 36966 35710 37018
rect 35722 36966 35774 37018
rect 35786 36966 35838 37018
rect 35850 36966 35902 37018
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 35594 35878 35646 35930
rect 35658 35878 35710 35930
rect 35722 35878 35774 35930
rect 35786 35878 35838 35930
rect 35850 35878 35902 35930
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 35594 34790 35646 34842
rect 35658 34790 35710 34842
rect 35722 34790 35774 34842
rect 35786 34790 35838 34842
rect 35850 34790 35902 34842
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 35594 33702 35646 33754
rect 35658 33702 35710 33754
rect 35722 33702 35774 33754
rect 35786 33702 35838 33754
rect 35850 33702 35902 33754
rect 38844 33464 38896 33516
rect 38292 33303 38344 33312
rect 38292 33269 38301 33303
rect 38301 33269 38335 33303
rect 38335 33269 38344 33303
rect 38292 33260 38344 33269
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 35594 32614 35646 32666
rect 35658 32614 35710 32666
rect 35722 32614 35774 32666
rect 35786 32614 35838 32666
rect 35850 32614 35902 32666
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 35594 31526 35646 31578
rect 35658 31526 35710 31578
rect 35722 31526 35774 31578
rect 35786 31526 35838 31578
rect 35850 31526 35902 31578
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 35594 30438 35646 30490
rect 35658 30438 35710 30490
rect 35722 30438 35774 30490
rect 35786 30438 35838 30490
rect 35850 30438 35902 30490
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 35594 29350 35646 29402
rect 35658 29350 35710 29402
rect 35722 29350 35774 29402
rect 35786 29350 35838 29402
rect 35850 29350 35902 29402
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 35594 28262 35646 28314
rect 35658 28262 35710 28314
rect 35722 28262 35774 28314
rect 35786 28262 35838 28314
rect 35850 28262 35902 28314
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 35594 27174 35646 27226
rect 35658 27174 35710 27226
rect 35722 27174 35774 27226
rect 35786 27174 35838 27226
rect 35850 27174 35902 27226
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 35594 26086 35646 26138
rect 35658 26086 35710 26138
rect 35722 26086 35774 26138
rect 35786 26086 35838 26138
rect 35850 26086 35902 26138
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 940 25168 992 25220
rect 19616 25100 19668 25152
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 35594 24998 35646 25050
rect 35658 24998 35710 25050
rect 35722 24998 35774 25050
rect 35786 24998 35838 25050
rect 35850 24998 35902 25050
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 35594 23910 35646 23962
rect 35658 23910 35710 23962
rect 35722 23910 35774 23962
rect 35786 23910 35838 23962
rect 35850 23910 35902 23962
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 35594 22822 35646 22874
rect 35658 22822 35710 22874
rect 35722 22822 35774 22874
rect 35786 22822 35838 22874
rect 35850 22822 35902 22874
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 35594 21734 35646 21786
rect 35658 21734 35710 21786
rect 35722 21734 35774 21786
rect 35786 21734 35838 21786
rect 35850 21734 35902 21786
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 35594 20646 35646 20698
rect 35658 20646 35710 20698
rect 35722 20646 35774 20698
rect 35786 20646 35838 20698
rect 35850 20646 35902 20698
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 35594 19558 35646 19610
rect 35658 19558 35710 19610
rect 35722 19558 35774 19610
rect 35786 19558 35838 19610
rect 35850 19558 35902 19610
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 35594 18470 35646 18522
rect 35658 18470 35710 18522
rect 35722 18470 35774 18522
rect 35786 18470 35838 18522
rect 35850 18470 35902 18522
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 35594 17382 35646 17434
rect 35658 17382 35710 17434
rect 35722 17382 35774 17434
rect 35786 17382 35838 17434
rect 35850 17382 35902 17434
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 35594 16294 35646 16346
rect 35658 16294 35710 16346
rect 35722 16294 35774 16346
rect 35786 16294 35838 16346
rect 35850 16294 35902 16346
rect 23664 16099 23716 16108
rect 23664 16065 23673 16099
rect 23673 16065 23707 16099
rect 23707 16065 23716 16099
rect 23664 16056 23716 16065
rect 33692 16056 33744 16108
rect 22376 15988 22428 16040
rect 24216 15988 24268 16040
rect 22284 15895 22336 15904
rect 22284 15861 22293 15895
rect 22293 15861 22327 15895
rect 22327 15861 22336 15895
rect 22284 15852 22336 15861
rect 23940 15895 23992 15904
rect 23940 15861 23949 15895
rect 23949 15861 23983 15895
rect 23983 15861 23992 15895
rect 23940 15852 23992 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 22284 15648 22336 15700
rect 23940 15648 23992 15700
rect 21088 15444 21140 15496
rect 20536 15351 20588 15360
rect 20536 15317 20545 15351
rect 20545 15317 20579 15351
rect 20579 15317 20588 15351
rect 20536 15308 20588 15317
rect 21180 15351 21232 15360
rect 21180 15317 21189 15351
rect 21189 15317 21223 15351
rect 21223 15317 21232 15351
rect 21180 15308 21232 15317
rect 21916 15444 21968 15496
rect 22284 15512 22336 15564
rect 22928 15444 22980 15496
rect 38292 15444 38344 15496
rect 22468 15351 22520 15360
rect 22468 15317 22477 15351
rect 22477 15317 22511 15351
rect 22511 15317 22520 15351
rect 22468 15308 22520 15317
rect 24952 15351 25004 15360
rect 24952 15317 24961 15351
rect 24961 15317 24995 15351
rect 24995 15317 25004 15351
rect 24952 15308 25004 15317
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 35594 15206 35646 15258
rect 35658 15206 35710 15258
rect 35722 15206 35774 15258
rect 35786 15206 35838 15258
rect 35850 15206 35902 15258
rect 20536 15104 20588 15156
rect 21088 15104 21140 15156
rect 22192 15147 22244 15156
rect 22192 15113 22201 15147
rect 22201 15113 22235 15147
rect 22235 15113 22244 15147
rect 22192 15104 22244 15113
rect 22468 15104 22520 15156
rect 23664 15147 23716 15156
rect 23664 15113 23673 15147
rect 23673 15113 23707 15147
rect 23707 15113 23716 15147
rect 23664 15104 23716 15113
rect 24952 15104 25004 15156
rect 18972 15011 19024 15020
rect 18972 14977 18981 15011
rect 18981 14977 19015 15011
rect 19015 14977 19024 15011
rect 18972 14968 19024 14977
rect 22284 14968 22336 15020
rect 18788 14807 18840 14816
rect 18788 14773 18797 14807
rect 18797 14773 18831 14807
rect 18831 14773 18840 14807
rect 18788 14764 18840 14773
rect 20536 14900 20588 14952
rect 21916 14900 21968 14952
rect 22928 14900 22980 14952
rect 24492 14968 24544 15020
rect 24032 14900 24084 14952
rect 25412 14968 25464 15020
rect 20720 14764 20772 14816
rect 22836 14764 22888 14816
rect 25044 14764 25096 14816
rect 25320 14807 25372 14816
rect 25320 14773 25329 14807
rect 25329 14773 25363 14807
rect 25363 14773 25372 14807
rect 25320 14764 25372 14773
rect 25504 14807 25556 14816
rect 25504 14773 25513 14807
rect 25513 14773 25547 14807
rect 25547 14773 25556 14807
rect 25504 14764 25556 14773
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 18972 14560 19024 14612
rect 20720 14560 20772 14612
rect 22376 14603 22428 14612
rect 22376 14569 22385 14603
rect 22385 14569 22419 14603
rect 22419 14569 22428 14603
rect 22376 14560 22428 14569
rect 20076 14424 20128 14476
rect 20536 14424 20588 14476
rect 25044 14492 25096 14544
rect 21916 14424 21968 14476
rect 22836 14424 22888 14476
rect 24032 14424 24084 14476
rect 26240 14424 26292 14476
rect 27160 14424 27212 14476
rect 27528 14424 27580 14476
rect 19616 14399 19668 14408
rect 19616 14365 19625 14399
rect 19625 14365 19659 14399
rect 19659 14365 19668 14399
rect 19616 14356 19668 14365
rect 22192 14356 22244 14408
rect 21180 14288 21232 14340
rect 25228 14356 25280 14408
rect 25320 14356 25372 14408
rect 19708 14263 19760 14272
rect 19708 14229 19717 14263
rect 19717 14229 19751 14263
rect 19751 14229 19760 14263
rect 19708 14220 19760 14229
rect 25412 14288 25464 14340
rect 27344 14288 27396 14340
rect 27896 14331 27948 14340
rect 27896 14297 27905 14331
rect 27905 14297 27939 14331
rect 27939 14297 27948 14331
rect 27896 14288 27948 14297
rect 22284 14220 22336 14272
rect 23664 14220 23716 14272
rect 24400 14263 24452 14272
rect 24400 14229 24409 14263
rect 24409 14229 24443 14263
rect 24443 14229 24452 14263
rect 24400 14220 24452 14229
rect 25780 14263 25832 14272
rect 25780 14229 25789 14263
rect 25789 14229 25823 14263
rect 25823 14229 25832 14263
rect 25780 14220 25832 14229
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 35594 14118 35646 14170
rect 35658 14118 35710 14170
rect 35722 14118 35774 14170
rect 35786 14118 35838 14170
rect 35850 14118 35902 14170
rect 19708 14016 19760 14068
rect 18788 13948 18840 14000
rect 20628 13948 20680 14000
rect 22284 14016 22336 14068
rect 21916 13948 21968 14000
rect 20904 13880 20956 13932
rect 23664 13948 23716 14000
rect 25504 14016 25556 14068
rect 25780 14016 25832 14068
rect 27896 14059 27948 14068
rect 27896 14025 27905 14059
rect 27905 14025 27939 14059
rect 27939 14025 27948 14059
rect 27896 14016 27948 14025
rect 26700 13948 26752 14000
rect 27712 13923 27764 13932
rect 27712 13889 27721 13923
rect 27721 13889 27755 13923
rect 27755 13889 27764 13923
rect 27712 13880 27764 13889
rect 18604 13855 18656 13864
rect 18604 13821 18613 13855
rect 18613 13821 18647 13855
rect 18647 13821 18656 13855
rect 18604 13812 18656 13821
rect 21916 13855 21968 13864
rect 21916 13821 21925 13855
rect 21925 13821 21959 13855
rect 21959 13821 21968 13855
rect 21916 13812 21968 13821
rect 23204 13855 23256 13864
rect 23204 13821 23213 13855
rect 23213 13821 23247 13855
rect 23247 13821 23256 13855
rect 23204 13812 23256 13821
rect 24492 13812 24544 13864
rect 24860 13855 24912 13864
rect 24860 13821 24869 13855
rect 24869 13821 24903 13855
rect 24903 13821 24912 13855
rect 24860 13812 24912 13821
rect 25872 13812 25924 13864
rect 22192 13676 22244 13728
rect 25228 13676 25280 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 10140 13472 10192 13524
rect 21916 13472 21968 13524
rect 23204 13515 23256 13524
rect 23204 13481 23213 13515
rect 23213 13481 23247 13515
rect 23247 13481 23256 13515
rect 23204 13472 23256 13481
rect 24032 13472 24084 13524
rect 19616 13336 19668 13388
rect 20904 13404 20956 13456
rect 27712 13472 27764 13524
rect 19432 13311 19484 13320
rect 19432 13277 19441 13311
rect 19441 13277 19475 13311
rect 19475 13277 19484 13311
rect 19432 13268 19484 13277
rect 19984 13132 20036 13184
rect 20720 13268 20772 13320
rect 22284 13268 22336 13320
rect 21180 13243 21232 13252
rect 21180 13209 21189 13243
rect 21189 13209 21223 13243
rect 21223 13209 21232 13243
rect 21180 13200 21232 13209
rect 22008 13132 22060 13184
rect 22928 13132 22980 13184
rect 24032 13379 24084 13388
rect 24032 13345 24041 13379
rect 24041 13345 24075 13379
rect 24075 13345 24084 13379
rect 24032 13336 24084 13345
rect 24216 13336 24268 13388
rect 24400 13336 24452 13388
rect 24860 13379 24912 13388
rect 24860 13345 24869 13379
rect 24869 13345 24903 13379
rect 24903 13345 24912 13379
rect 24860 13336 24912 13345
rect 25320 13268 25372 13320
rect 27528 13268 27580 13320
rect 28080 13311 28132 13320
rect 26240 13200 26292 13252
rect 27160 13243 27212 13252
rect 27160 13209 27169 13243
rect 27169 13209 27203 13243
rect 27203 13209 27212 13243
rect 27160 13200 27212 13209
rect 26608 13132 26660 13184
rect 28080 13277 28089 13311
rect 28089 13277 28123 13311
rect 28123 13277 28132 13311
rect 28080 13268 28132 13277
rect 29920 13132 29972 13184
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 35594 13030 35646 13082
rect 35658 13030 35710 13082
rect 35722 13030 35774 13082
rect 35786 13030 35838 13082
rect 35850 13030 35902 13082
rect 21180 12928 21232 12980
rect 22192 12928 22244 12980
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 19984 12860 20036 12912
rect 21456 12835 21508 12844
rect 21456 12801 21465 12835
rect 21465 12801 21499 12835
rect 21499 12801 21508 12835
rect 21456 12792 21508 12801
rect 22836 12835 22888 12844
rect 22836 12801 22870 12835
rect 22870 12801 22888 12835
rect 22836 12792 22888 12801
rect 20076 12767 20128 12776
rect 20076 12733 20085 12767
rect 20085 12733 20119 12767
rect 20119 12733 20128 12767
rect 20076 12724 20128 12733
rect 21088 12767 21140 12776
rect 21088 12733 21097 12767
rect 21097 12733 21131 12767
rect 21131 12733 21140 12767
rect 21088 12724 21140 12733
rect 19524 12588 19576 12640
rect 22376 12724 22428 12776
rect 23204 12724 23256 12776
rect 26240 12928 26292 12980
rect 27344 12928 27396 12980
rect 24400 12835 24452 12844
rect 24400 12801 24409 12835
rect 24409 12801 24443 12835
rect 24443 12801 24452 12835
rect 24400 12792 24452 12801
rect 25228 12792 25280 12844
rect 22560 12656 22612 12708
rect 24676 12767 24728 12776
rect 24676 12733 24685 12767
rect 24685 12733 24719 12767
rect 24719 12733 24728 12767
rect 24676 12724 24728 12733
rect 25044 12724 25096 12776
rect 25964 12724 26016 12776
rect 22928 12588 22980 12640
rect 23664 12631 23716 12640
rect 23664 12597 23673 12631
rect 23673 12597 23707 12631
rect 23707 12597 23716 12631
rect 23664 12588 23716 12597
rect 23756 12631 23808 12640
rect 23756 12597 23765 12631
rect 23765 12597 23799 12631
rect 23799 12597 23808 12631
rect 23756 12588 23808 12597
rect 24952 12699 25004 12708
rect 24952 12665 24961 12699
rect 24961 12665 24995 12699
rect 24995 12665 25004 12699
rect 24952 12656 25004 12665
rect 25504 12656 25556 12708
rect 26240 12767 26292 12776
rect 26240 12733 26249 12767
rect 26249 12733 26283 12767
rect 26283 12733 26292 12767
rect 26240 12724 26292 12733
rect 26792 12835 26844 12844
rect 26792 12801 26801 12835
rect 26801 12801 26835 12835
rect 26835 12801 26844 12835
rect 26792 12792 26844 12801
rect 28816 12792 28868 12844
rect 26424 12724 26476 12776
rect 26332 12656 26384 12708
rect 27712 12767 27764 12776
rect 27712 12733 27721 12767
rect 27721 12733 27755 12767
rect 27755 12733 27764 12767
rect 27712 12724 27764 12733
rect 29552 12724 29604 12776
rect 24400 12588 24452 12640
rect 24492 12588 24544 12640
rect 27528 12588 27580 12640
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 18604 12248 18656 12300
rect 19984 12384 20036 12436
rect 20812 12248 20864 12300
rect 21088 12384 21140 12436
rect 21456 12384 21508 12436
rect 23664 12384 23716 12436
rect 27712 12384 27764 12436
rect 22928 12291 22980 12300
rect 22928 12257 22937 12291
rect 22937 12257 22971 12291
rect 22971 12257 22980 12291
rect 22928 12248 22980 12257
rect 18236 12087 18288 12096
rect 18236 12053 18245 12087
rect 18245 12053 18279 12087
rect 18279 12053 18288 12087
rect 18236 12044 18288 12053
rect 20628 12180 20680 12232
rect 22008 12180 22060 12232
rect 23848 12223 23900 12232
rect 23848 12189 23857 12223
rect 23857 12189 23891 12223
rect 23891 12189 23900 12223
rect 23848 12180 23900 12189
rect 19432 12112 19484 12164
rect 19524 12155 19576 12164
rect 19524 12121 19533 12155
rect 19533 12121 19567 12155
rect 19567 12121 19576 12155
rect 19524 12112 19576 12121
rect 25412 12223 25464 12232
rect 25412 12189 25421 12223
rect 25421 12189 25455 12223
rect 25455 12189 25464 12223
rect 25412 12180 25464 12189
rect 25872 12291 25924 12300
rect 25872 12257 25881 12291
rect 25881 12257 25915 12291
rect 25915 12257 25924 12291
rect 25872 12248 25924 12257
rect 26424 12316 26476 12368
rect 26608 12291 26660 12300
rect 26608 12257 26617 12291
rect 26617 12257 26651 12291
rect 26651 12257 26660 12291
rect 26608 12248 26660 12257
rect 29552 12316 29604 12368
rect 25964 12180 26016 12232
rect 26240 12223 26292 12232
rect 26240 12189 26249 12223
rect 26249 12189 26283 12223
rect 26283 12189 26292 12223
rect 26240 12180 26292 12189
rect 26884 12223 26936 12232
rect 26884 12189 26893 12223
rect 26893 12189 26927 12223
rect 26927 12189 26936 12223
rect 26884 12180 26936 12189
rect 26976 12180 27028 12232
rect 28080 12248 28132 12300
rect 27252 12223 27304 12232
rect 27252 12189 27261 12223
rect 27261 12189 27295 12223
rect 27295 12189 27304 12223
rect 27252 12180 27304 12189
rect 18696 12087 18748 12096
rect 18696 12053 18705 12087
rect 18705 12053 18739 12087
rect 18739 12053 18748 12087
rect 18696 12044 18748 12053
rect 18788 12087 18840 12096
rect 18788 12053 18797 12087
rect 18797 12053 18831 12087
rect 18831 12053 18840 12087
rect 18788 12044 18840 12053
rect 24584 12044 24636 12096
rect 26424 12112 26476 12164
rect 28172 12223 28224 12232
rect 28172 12189 28181 12223
rect 28181 12189 28215 12223
rect 28215 12189 28224 12223
rect 28172 12180 28224 12189
rect 28724 12180 28776 12232
rect 25228 12087 25280 12096
rect 25228 12053 25237 12087
rect 25237 12053 25271 12087
rect 25271 12053 25280 12087
rect 25228 12044 25280 12053
rect 25964 12087 26016 12096
rect 25964 12053 25973 12087
rect 25973 12053 26007 12087
rect 26007 12053 26016 12087
rect 25964 12044 26016 12053
rect 27620 12087 27672 12096
rect 27620 12053 27629 12087
rect 27629 12053 27663 12087
rect 27663 12053 27672 12087
rect 27620 12044 27672 12053
rect 29736 12044 29788 12096
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 35594 11942 35646 11994
rect 35658 11942 35710 11994
rect 35722 11942 35774 11994
rect 35786 11942 35838 11994
rect 35850 11942 35902 11994
rect 18236 11840 18288 11892
rect 18604 11840 18656 11892
rect 20444 11883 20496 11892
rect 20444 11849 20453 11883
rect 20453 11849 20487 11883
rect 20487 11849 20496 11883
rect 20444 11840 20496 11849
rect 26424 11840 26476 11892
rect 28172 11840 28224 11892
rect 20628 11772 20680 11824
rect 22100 11772 22152 11824
rect 22192 11747 22244 11756
rect 22192 11713 22201 11747
rect 22201 11713 22235 11747
rect 22235 11713 22244 11747
rect 22192 11704 22244 11713
rect 23204 11772 23256 11824
rect 23572 11772 23624 11824
rect 24676 11772 24728 11824
rect 22560 11636 22612 11688
rect 25136 11704 25188 11756
rect 26332 11747 26384 11756
rect 22928 11636 22980 11688
rect 20812 11568 20864 11620
rect 23756 11636 23808 11688
rect 26332 11713 26341 11747
rect 26341 11713 26375 11747
rect 26375 11713 26384 11747
rect 26332 11704 26384 11713
rect 26884 11704 26936 11756
rect 28816 11704 28868 11756
rect 29644 11747 29696 11756
rect 29644 11713 29653 11747
rect 29653 11713 29687 11747
rect 29687 11713 29696 11747
rect 29644 11704 29696 11713
rect 21824 11543 21876 11552
rect 21824 11509 21833 11543
rect 21833 11509 21867 11543
rect 21867 11509 21876 11543
rect 21824 11500 21876 11509
rect 23112 11500 23164 11552
rect 24584 11500 24636 11552
rect 25596 11568 25648 11620
rect 27528 11679 27580 11688
rect 27528 11645 27537 11679
rect 27537 11645 27571 11679
rect 27571 11645 27580 11679
rect 27528 11636 27580 11645
rect 27804 11679 27856 11688
rect 27804 11645 27813 11679
rect 27813 11645 27847 11679
rect 27847 11645 27856 11679
rect 27804 11636 27856 11645
rect 29920 11568 29972 11620
rect 38200 11568 38252 11620
rect 24860 11543 24912 11552
rect 24860 11509 24869 11543
rect 24869 11509 24903 11543
rect 24903 11509 24912 11543
rect 24860 11500 24912 11509
rect 25044 11500 25096 11552
rect 26424 11500 26476 11552
rect 26608 11500 26660 11552
rect 27620 11500 27672 11552
rect 29736 11500 29788 11552
rect 29828 11543 29880 11552
rect 29828 11509 29837 11543
rect 29837 11509 29871 11543
rect 29871 11509 29880 11543
rect 29828 11500 29880 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 18788 11296 18840 11348
rect 20812 11296 20864 11348
rect 22100 11296 22152 11348
rect 23020 11296 23072 11348
rect 25228 11296 25280 11348
rect 25320 11296 25372 11348
rect 25964 11296 26016 11348
rect 26148 11296 26200 11348
rect 26884 11296 26936 11348
rect 27804 11339 27856 11348
rect 27804 11305 27813 11339
rect 27813 11305 27847 11339
rect 27847 11305 27856 11339
rect 27804 11296 27856 11305
rect 27896 11339 27948 11348
rect 27896 11305 27905 11339
rect 27905 11305 27939 11339
rect 27939 11305 27948 11339
rect 27896 11296 27948 11305
rect 29552 11296 29604 11348
rect 29828 11296 29880 11348
rect 20444 11160 20496 11212
rect 23204 11228 23256 11280
rect 23572 11228 23624 11280
rect 22192 11160 22244 11212
rect 20628 11092 20680 11144
rect 20996 11067 21048 11076
rect 20996 11033 21005 11067
rect 21005 11033 21039 11067
rect 21039 11033 21048 11067
rect 20996 11024 21048 11033
rect 22928 11024 22980 11076
rect 22836 10999 22888 11008
rect 22836 10965 22845 10999
rect 22845 10965 22879 10999
rect 22879 10965 22888 10999
rect 22836 10956 22888 10965
rect 23848 11092 23900 11144
rect 25136 11203 25188 11212
rect 25136 11169 25145 11203
rect 25145 11169 25179 11203
rect 25179 11169 25188 11203
rect 25136 11160 25188 11169
rect 24400 11092 24452 11144
rect 24952 11092 25004 11144
rect 25044 11135 25096 11144
rect 25044 11101 25053 11135
rect 25053 11101 25087 11135
rect 25087 11101 25096 11135
rect 25044 11092 25096 11101
rect 25412 11092 25464 11144
rect 26608 11228 26660 11280
rect 26516 11203 26568 11212
rect 26516 11169 26525 11203
rect 26525 11169 26559 11203
rect 26559 11169 26568 11203
rect 26516 11160 26568 11169
rect 27344 11228 27396 11280
rect 23204 11067 23256 11076
rect 23204 11033 23213 11067
rect 23213 11033 23247 11067
rect 23247 11033 23256 11067
rect 23204 11024 23256 11033
rect 25320 11024 25372 11076
rect 25596 11024 25648 11076
rect 25872 11024 25924 11076
rect 26976 11092 27028 11144
rect 27620 11135 27672 11144
rect 27620 11101 27629 11135
rect 27629 11101 27663 11135
rect 27663 11101 27672 11135
rect 27620 11092 27672 11101
rect 27804 11092 27856 11144
rect 29920 11160 29972 11212
rect 27252 11067 27304 11076
rect 27252 11033 27261 11067
rect 27261 11033 27295 11067
rect 27295 11033 27304 11067
rect 29552 11135 29604 11144
rect 29552 11101 29561 11135
rect 29561 11101 29595 11135
rect 29595 11101 29604 11135
rect 29552 11092 29604 11101
rect 29644 11135 29696 11144
rect 29644 11101 29653 11135
rect 29653 11101 29687 11135
rect 29687 11101 29696 11135
rect 29644 11092 29696 11101
rect 29736 11092 29788 11144
rect 27252 11024 27304 11033
rect 23480 10956 23532 11008
rect 23940 10956 23992 11008
rect 24676 10956 24728 11008
rect 26424 10999 26476 11008
rect 26424 10965 26433 10999
rect 26433 10965 26467 10999
rect 26467 10965 26476 10999
rect 26424 10956 26476 10965
rect 26700 10999 26752 11008
rect 26700 10965 26709 10999
rect 26709 10965 26743 10999
rect 26743 10965 26752 10999
rect 26700 10956 26752 10965
rect 26884 10956 26936 11008
rect 27344 10956 27396 11008
rect 30012 10999 30064 11008
rect 30012 10965 30021 10999
rect 30021 10965 30055 10999
rect 30055 10965 30064 10999
rect 30012 10956 30064 10965
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 35594 10854 35646 10906
rect 35658 10854 35710 10906
rect 35722 10854 35774 10906
rect 35786 10854 35838 10906
rect 35850 10854 35902 10906
rect 20996 10752 21048 10804
rect 21824 10752 21876 10804
rect 20812 10616 20864 10668
rect 22836 10752 22888 10804
rect 23572 10795 23624 10804
rect 23572 10761 23581 10795
rect 23581 10761 23615 10795
rect 23615 10761 23624 10795
rect 23572 10752 23624 10761
rect 23756 10795 23808 10804
rect 23756 10761 23765 10795
rect 23765 10761 23799 10795
rect 23799 10761 23808 10795
rect 23756 10752 23808 10761
rect 23848 10752 23900 10804
rect 25228 10752 25280 10804
rect 26332 10752 26384 10804
rect 26424 10752 26476 10804
rect 26976 10752 27028 10804
rect 27344 10795 27396 10804
rect 27344 10761 27353 10795
rect 27353 10761 27387 10795
rect 27387 10761 27396 10795
rect 27344 10752 27396 10761
rect 27804 10752 27856 10804
rect 27896 10752 27948 10804
rect 29644 10752 29696 10804
rect 23388 10684 23440 10736
rect 23940 10659 23992 10668
rect 23940 10625 23949 10659
rect 23949 10625 23983 10659
rect 23983 10625 23992 10659
rect 23940 10616 23992 10625
rect 26240 10727 26292 10736
rect 26240 10693 26249 10727
rect 26249 10693 26283 10727
rect 26283 10693 26292 10727
rect 26240 10684 26292 10693
rect 24860 10616 24912 10668
rect 25872 10616 25924 10668
rect 27252 10684 27304 10736
rect 28816 10684 28868 10736
rect 25688 10548 25740 10600
rect 24676 10480 24728 10532
rect 27620 10548 27672 10600
rect 22468 10412 22520 10464
rect 25964 10412 26016 10464
rect 26700 10412 26752 10464
rect 27160 10412 27212 10464
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 20812 10208 20864 10260
rect 23480 10251 23532 10260
rect 23480 10217 23489 10251
rect 23489 10217 23523 10251
rect 23523 10217 23532 10251
rect 23480 10208 23532 10217
rect 24400 10072 24452 10124
rect 24492 10115 24544 10124
rect 24492 10081 24501 10115
rect 24501 10081 24535 10115
rect 24535 10081 24544 10115
rect 24492 10072 24544 10081
rect 24584 10115 24636 10124
rect 24584 10081 24593 10115
rect 24593 10081 24627 10115
rect 24627 10081 24636 10115
rect 24584 10072 24636 10081
rect 23296 10047 23348 10056
rect 23296 10013 23305 10047
rect 23305 10013 23339 10047
rect 23339 10013 23348 10047
rect 23296 10004 23348 10013
rect 22468 9936 22520 9988
rect 22928 9936 22980 9988
rect 24952 10072 25004 10124
rect 25136 10208 25188 10260
rect 25136 10072 25188 10124
rect 25504 10208 25556 10260
rect 27528 10251 27580 10260
rect 27528 10217 27537 10251
rect 27537 10217 27571 10251
rect 27571 10217 27580 10251
rect 27528 10208 27580 10217
rect 25412 10004 25464 10056
rect 25780 10047 25832 10056
rect 25780 10013 25789 10047
rect 25789 10013 25823 10047
rect 25823 10013 25832 10047
rect 25780 10004 25832 10013
rect 25964 10004 26016 10056
rect 26240 10004 26292 10056
rect 28080 10047 28132 10056
rect 28080 10013 28089 10047
rect 28089 10013 28123 10047
rect 28123 10013 28132 10047
rect 28080 10004 28132 10013
rect 30012 10004 30064 10056
rect 30104 10047 30156 10056
rect 30104 10013 30113 10047
rect 30113 10013 30147 10047
rect 30147 10013 30156 10047
rect 30104 10004 30156 10013
rect 27252 9936 27304 9988
rect 22744 9911 22796 9920
rect 22744 9877 22753 9911
rect 22753 9877 22787 9911
rect 22787 9877 22796 9911
rect 22744 9868 22796 9877
rect 24952 9911 25004 9920
rect 24952 9877 24961 9911
rect 24961 9877 24995 9911
rect 24995 9877 25004 9911
rect 24952 9868 25004 9877
rect 25504 9868 25556 9920
rect 25596 9868 25648 9920
rect 25964 9911 26016 9920
rect 25964 9877 25973 9911
rect 25973 9877 26007 9911
rect 26007 9877 26016 9911
rect 25964 9868 26016 9877
rect 27712 9868 27764 9920
rect 28172 9979 28224 9988
rect 28172 9945 28181 9979
rect 28181 9945 28215 9979
rect 28215 9945 28224 9979
rect 28172 9936 28224 9945
rect 28632 9936 28684 9988
rect 28724 9979 28776 9988
rect 28724 9945 28733 9979
rect 28733 9945 28767 9979
rect 28767 9945 28776 9979
rect 28724 9936 28776 9945
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 35594 9766 35646 9818
rect 35658 9766 35710 9818
rect 35722 9766 35774 9818
rect 35786 9766 35838 9818
rect 35850 9766 35902 9818
rect 23020 9596 23072 9648
rect 24952 9664 25004 9716
rect 24584 9596 24636 9648
rect 25044 9596 25096 9648
rect 22744 9528 22796 9580
rect 25504 9639 25556 9648
rect 25504 9605 25513 9639
rect 25513 9605 25547 9639
rect 25547 9605 25556 9639
rect 25504 9596 25556 9605
rect 25688 9707 25740 9716
rect 25688 9673 25697 9707
rect 25697 9673 25731 9707
rect 25731 9673 25740 9707
rect 25688 9664 25740 9673
rect 25872 9707 25924 9716
rect 25872 9673 25881 9707
rect 25881 9673 25915 9707
rect 25915 9673 25924 9707
rect 25872 9664 25924 9673
rect 26148 9664 26200 9716
rect 26240 9664 26292 9716
rect 30104 9664 30156 9716
rect 24308 9503 24360 9512
rect 24308 9469 24317 9503
rect 24317 9469 24351 9503
rect 24351 9469 24360 9503
rect 24308 9460 24360 9469
rect 24676 9460 24728 9512
rect 25872 9528 25924 9580
rect 26148 9571 26200 9580
rect 26148 9537 26157 9571
rect 26157 9537 26191 9571
rect 26191 9537 26200 9571
rect 26148 9528 26200 9537
rect 25964 9460 26016 9512
rect 25504 9392 25556 9444
rect 21732 9324 21784 9376
rect 22836 9367 22888 9376
rect 22836 9333 22845 9367
rect 22845 9333 22879 9367
rect 22879 9333 22888 9367
rect 22836 9324 22888 9333
rect 24676 9367 24728 9376
rect 24676 9333 24685 9367
rect 24685 9333 24719 9367
rect 24719 9333 24728 9367
rect 24676 9324 24728 9333
rect 25228 9324 25280 9376
rect 25320 9367 25372 9376
rect 25320 9333 25329 9367
rect 25329 9333 25363 9367
rect 25363 9333 25372 9367
rect 25320 9324 25372 9333
rect 25412 9324 25464 9376
rect 26608 9571 26660 9580
rect 26608 9537 26617 9571
rect 26617 9537 26651 9571
rect 26651 9537 26660 9571
rect 26608 9528 26660 9537
rect 27252 9596 27304 9648
rect 27712 9639 27764 9648
rect 27712 9605 27721 9639
rect 27721 9605 27755 9639
rect 27755 9605 27764 9639
rect 27712 9596 27764 9605
rect 28264 9596 28316 9648
rect 26700 9460 26752 9512
rect 26884 9460 26936 9512
rect 27068 9503 27120 9512
rect 27068 9469 27077 9503
rect 27077 9469 27111 9503
rect 27111 9469 27120 9503
rect 27068 9460 27120 9469
rect 27436 9503 27488 9512
rect 27436 9469 27445 9503
rect 27445 9469 27479 9503
rect 27479 9469 27488 9503
rect 27436 9460 27488 9469
rect 27344 9435 27396 9444
rect 27344 9401 27353 9435
rect 27353 9401 27387 9435
rect 27387 9401 27396 9435
rect 27344 9392 27396 9401
rect 26516 9324 26568 9376
rect 26976 9324 27028 9376
rect 27160 9367 27212 9376
rect 27160 9333 27169 9367
rect 27169 9333 27203 9367
rect 27203 9333 27212 9367
rect 27160 9324 27212 9333
rect 28448 9324 28500 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 23296 9120 23348 9172
rect 24308 9120 24360 9172
rect 24584 9120 24636 9172
rect 24676 9120 24728 9172
rect 25780 9120 25832 9172
rect 26792 9120 26844 9172
rect 21824 8984 21876 9036
rect 22836 8984 22888 9036
rect 23020 8984 23072 9036
rect 22560 8916 22612 8968
rect 22928 8916 22980 8968
rect 25504 8984 25556 9036
rect 26700 9052 26752 9104
rect 28264 9120 28316 9172
rect 28540 9163 28592 9172
rect 28540 9129 28549 9163
rect 28549 9129 28583 9163
rect 28583 9129 28592 9163
rect 28540 9120 28592 9129
rect 28632 9120 28684 9172
rect 30012 9120 30064 9172
rect 21456 8891 21508 8900
rect 21456 8857 21465 8891
rect 21465 8857 21499 8891
rect 21499 8857 21508 8891
rect 21456 8848 21508 8857
rect 25780 8848 25832 8900
rect 27344 8984 27396 9036
rect 29736 9052 29788 9104
rect 28080 8984 28132 9036
rect 25596 8780 25648 8832
rect 26148 8780 26200 8832
rect 28172 8916 28224 8968
rect 27068 8780 27120 8832
rect 28724 8848 28776 8900
rect 27804 8780 27856 8832
rect 27896 8823 27948 8832
rect 27896 8789 27905 8823
rect 27905 8789 27939 8823
rect 27939 8789 27948 8823
rect 27896 8780 27948 8789
rect 28080 8823 28132 8832
rect 28080 8789 28089 8823
rect 28089 8789 28123 8823
rect 28123 8789 28132 8823
rect 28080 8780 28132 8789
rect 29552 8780 29604 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 35594 8678 35646 8730
rect 35658 8678 35710 8730
rect 35722 8678 35774 8730
rect 35786 8678 35838 8730
rect 35850 8678 35902 8730
rect 21456 8619 21508 8628
rect 21456 8585 21465 8619
rect 21465 8585 21499 8619
rect 21499 8585 21508 8619
rect 21456 8576 21508 8585
rect 21732 8576 21784 8628
rect 22560 8508 22612 8560
rect 21824 8483 21876 8492
rect 21824 8449 21833 8483
rect 21833 8449 21867 8483
rect 21867 8449 21876 8483
rect 21824 8440 21876 8449
rect 25780 8508 25832 8560
rect 27436 8576 27488 8628
rect 28908 8576 28960 8628
rect 22100 8415 22152 8424
rect 22100 8381 22109 8415
rect 22109 8381 22143 8415
rect 22143 8381 22152 8415
rect 22100 8372 22152 8381
rect 23572 8279 23624 8288
rect 23572 8245 23581 8279
rect 23581 8245 23615 8279
rect 23615 8245 23624 8279
rect 23572 8236 23624 8245
rect 23664 8279 23716 8288
rect 23664 8245 23673 8279
rect 23673 8245 23707 8279
rect 23707 8245 23716 8279
rect 23664 8236 23716 8245
rect 24032 8415 24084 8424
rect 24032 8381 24041 8415
rect 24041 8381 24075 8415
rect 24075 8381 24084 8415
rect 24032 8372 24084 8381
rect 26332 8483 26384 8492
rect 26332 8449 26341 8483
rect 26341 8449 26375 8483
rect 26375 8449 26384 8483
rect 26332 8440 26384 8449
rect 26424 8483 26476 8492
rect 26424 8449 26459 8483
rect 26459 8449 26476 8483
rect 27896 8508 27948 8560
rect 28264 8508 28316 8560
rect 29644 8551 29696 8560
rect 29644 8517 29653 8551
rect 29653 8517 29687 8551
rect 29687 8517 29696 8551
rect 29644 8508 29696 8517
rect 26424 8440 26476 8449
rect 27528 8440 27580 8492
rect 27620 8483 27672 8492
rect 27620 8449 27629 8483
rect 27629 8449 27663 8483
rect 27663 8449 27672 8483
rect 27620 8440 27672 8449
rect 27804 8483 27856 8492
rect 27804 8449 27813 8483
rect 27813 8449 27847 8483
rect 27847 8449 27856 8483
rect 27804 8440 27856 8449
rect 28080 8440 28132 8492
rect 38200 8576 38252 8628
rect 26884 8304 26936 8356
rect 24492 8236 24544 8288
rect 30012 8440 30064 8492
rect 30196 8483 30248 8492
rect 30196 8449 30205 8483
rect 30205 8449 30239 8483
rect 30239 8449 30248 8483
rect 30196 8440 30248 8449
rect 28632 8372 28684 8424
rect 30564 8483 30616 8492
rect 30564 8449 30573 8483
rect 30573 8449 30607 8483
rect 30607 8449 30616 8483
rect 30564 8440 30616 8449
rect 38844 8304 38896 8356
rect 28356 8236 28408 8288
rect 28448 8236 28500 8288
rect 29828 8236 29880 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 20812 8032 20864 8084
rect 21824 8032 21876 8084
rect 22100 8032 22152 8084
rect 23296 8032 23348 8084
rect 23664 8032 23716 8084
rect 24032 8032 24084 8084
rect 27068 8032 27120 8084
rect 27436 8032 27488 8084
rect 27988 8032 28040 8084
rect 28264 8032 28316 8084
rect 29276 8032 29328 8084
rect 29644 8032 29696 8084
rect 30564 8032 30616 8084
rect 22468 7828 22520 7880
rect 23572 7939 23624 7948
rect 23572 7905 23581 7939
rect 23581 7905 23615 7939
rect 23615 7905 23624 7939
rect 23572 7896 23624 7905
rect 23020 7828 23072 7880
rect 27804 7896 27856 7948
rect 26056 7871 26108 7880
rect 26056 7837 26065 7871
rect 26065 7837 26099 7871
rect 26099 7837 26108 7871
rect 26056 7828 26108 7837
rect 28632 7896 28684 7948
rect 29552 7939 29604 7948
rect 29552 7905 29561 7939
rect 29561 7905 29595 7939
rect 29595 7905 29604 7939
rect 29552 7896 29604 7905
rect 29736 7896 29788 7948
rect 22928 7803 22980 7812
rect 22928 7769 22937 7803
rect 22937 7769 22971 7803
rect 22971 7769 22980 7803
rect 22928 7760 22980 7769
rect 24492 7760 24544 7812
rect 25412 7692 25464 7744
rect 27896 7760 27948 7812
rect 28356 7871 28408 7880
rect 28356 7837 28365 7871
rect 28365 7837 28399 7871
rect 28399 7837 28408 7871
rect 28356 7828 28408 7837
rect 30012 7871 30064 7880
rect 30012 7837 30021 7871
rect 30021 7837 30055 7871
rect 30055 7837 30064 7871
rect 30012 7828 30064 7837
rect 30288 7871 30340 7880
rect 30288 7837 30297 7871
rect 30297 7837 30331 7871
rect 30331 7837 30340 7871
rect 30288 7828 30340 7837
rect 26332 7692 26384 7744
rect 28448 7692 28500 7744
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 35594 7590 35646 7642
rect 35658 7590 35710 7642
rect 35722 7590 35774 7642
rect 35786 7590 35838 7642
rect 35850 7590 35902 7642
rect 22928 7488 22980 7540
rect 25872 7488 25924 7540
rect 30196 7488 30248 7540
rect 30288 7531 30340 7540
rect 30288 7497 30297 7531
rect 30297 7497 30331 7531
rect 30331 7497 30340 7531
rect 30288 7488 30340 7497
rect 22744 7327 22796 7336
rect 22744 7293 22753 7327
rect 22753 7293 22787 7327
rect 22787 7293 22796 7327
rect 22744 7284 22796 7293
rect 23020 7284 23072 7336
rect 23848 7395 23900 7404
rect 23848 7361 23857 7395
rect 23857 7361 23891 7395
rect 23891 7361 23900 7395
rect 23848 7352 23900 7361
rect 24492 7420 24544 7472
rect 24400 7395 24452 7404
rect 24400 7361 24409 7395
rect 24409 7361 24443 7395
rect 24443 7361 24452 7395
rect 24400 7352 24452 7361
rect 24860 7352 24912 7404
rect 26516 7395 26568 7404
rect 26516 7361 26525 7395
rect 26525 7361 26559 7395
rect 26559 7361 26568 7395
rect 26516 7352 26568 7361
rect 26608 7395 26660 7404
rect 26608 7361 26617 7395
rect 26617 7361 26651 7395
rect 26651 7361 26660 7395
rect 26608 7352 26660 7361
rect 26976 7352 27028 7404
rect 27896 7420 27948 7472
rect 27620 7352 27672 7404
rect 23664 7327 23716 7336
rect 23664 7293 23673 7327
rect 23673 7293 23707 7327
rect 23707 7293 23716 7327
rect 23664 7284 23716 7293
rect 27160 7327 27212 7336
rect 27160 7293 27169 7327
rect 27169 7293 27203 7327
rect 27203 7293 27212 7327
rect 27160 7284 27212 7293
rect 27344 7327 27396 7336
rect 27344 7293 27353 7327
rect 27353 7293 27387 7327
rect 27387 7293 27396 7327
rect 27344 7284 27396 7293
rect 27804 7327 27856 7336
rect 27804 7293 27813 7327
rect 27813 7293 27847 7327
rect 27847 7293 27856 7327
rect 27804 7284 27856 7293
rect 27896 7327 27948 7336
rect 27896 7293 27905 7327
rect 27905 7293 27939 7327
rect 27939 7293 27948 7327
rect 27896 7284 27948 7293
rect 28264 7395 28316 7404
rect 28264 7361 28273 7395
rect 28273 7361 28307 7395
rect 28307 7361 28316 7395
rect 28264 7352 28316 7361
rect 28448 7395 28500 7404
rect 28448 7361 28457 7395
rect 28457 7361 28491 7395
rect 28491 7361 28500 7395
rect 28448 7352 28500 7361
rect 28908 7420 28960 7472
rect 29092 7420 29144 7472
rect 29276 7420 29328 7472
rect 29828 7352 29880 7404
rect 20536 7191 20588 7200
rect 20536 7157 20545 7191
rect 20545 7157 20579 7191
rect 20579 7157 20588 7191
rect 20536 7148 20588 7157
rect 21824 7191 21876 7200
rect 21824 7157 21833 7191
rect 21833 7157 21867 7191
rect 21867 7157 21876 7191
rect 21824 7148 21876 7157
rect 27528 7216 27580 7268
rect 24124 7191 24176 7200
rect 24124 7157 24133 7191
rect 24133 7157 24167 7191
rect 24167 7157 24176 7191
rect 24124 7148 24176 7157
rect 24308 7148 24360 7200
rect 26700 7191 26752 7200
rect 26700 7157 26709 7191
rect 26709 7157 26743 7191
rect 26743 7157 26752 7191
rect 26700 7148 26752 7157
rect 27344 7148 27396 7200
rect 28356 7216 28408 7268
rect 28908 7148 28960 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 20536 6944 20588 6996
rect 24860 6987 24912 6996
rect 24860 6953 24869 6987
rect 24869 6953 24903 6987
rect 24903 6953 24912 6987
rect 24860 6944 24912 6953
rect 20812 6808 20864 6860
rect 22744 6808 22796 6860
rect 22192 6740 22244 6792
rect 22560 6740 22612 6792
rect 23480 6808 23532 6860
rect 23664 6851 23716 6860
rect 23664 6817 23673 6851
rect 23673 6817 23707 6851
rect 23707 6817 23716 6851
rect 23664 6808 23716 6817
rect 23848 6808 23900 6860
rect 24124 6740 24176 6792
rect 24400 6740 24452 6792
rect 24492 6740 24544 6792
rect 25504 6740 25556 6792
rect 26700 6944 26752 6996
rect 27804 6944 27856 6996
rect 28632 6987 28684 6996
rect 28632 6953 28641 6987
rect 28641 6953 28675 6987
rect 28675 6953 28684 6987
rect 28632 6944 28684 6953
rect 28816 6944 28868 6996
rect 29736 6944 29788 6996
rect 30012 6944 30064 6996
rect 26332 6876 26384 6928
rect 27160 6876 27212 6928
rect 26056 6783 26108 6792
rect 26056 6749 26065 6783
rect 26065 6749 26099 6783
rect 26099 6749 26108 6783
rect 26056 6740 26108 6749
rect 26332 6783 26384 6792
rect 26332 6749 26341 6783
rect 26341 6749 26375 6783
rect 26375 6749 26384 6783
rect 26332 6740 26384 6749
rect 22100 6715 22152 6724
rect 22100 6681 22109 6715
rect 22109 6681 22143 6715
rect 22143 6681 22152 6715
rect 22100 6672 22152 6681
rect 23112 6672 23164 6724
rect 20720 6604 20772 6656
rect 21824 6604 21876 6656
rect 23664 6604 23716 6656
rect 24400 6647 24452 6656
rect 24400 6613 24409 6647
rect 24409 6613 24443 6647
rect 24443 6613 24452 6647
rect 24400 6604 24452 6613
rect 25688 6647 25740 6656
rect 25688 6613 25697 6647
rect 25697 6613 25731 6647
rect 25731 6613 25740 6647
rect 25688 6604 25740 6613
rect 26608 6783 26660 6792
rect 26608 6749 26617 6783
rect 26617 6749 26651 6783
rect 26651 6749 26660 6783
rect 26608 6740 26660 6749
rect 26976 6740 27028 6792
rect 28908 6808 28960 6860
rect 26516 6672 26568 6724
rect 27436 6740 27488 6792
rect 27620 6740 27672 6792
rect 27712 6740 27764 6792
rect 28448 6740 28500 6792
rect 26056 6604 26108 6656
rect 26976 6604 27028 6656
rect 27436 6604 27488 6656
rect 28908 6672 28960 6724
rect 28356 6604 28408 6656
rect 28448 6647 28500 6656
rect 28448 6613 28457 6647
rect 28457 6613 28491 6647
rect 28491 6613 28500 6647
rect 28448 6604 28500 6613
rect 28816 6604 28868 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 35594 6502 35646 6554
rect 35658 6502 35710 6554
rect 35722 6502 35774 6554
rect 35786 6502 35838 6554
rect 35850 6502 35902 6554
rect 20812 6400 20864 6452
rect 23020 6400 23072 6452
rect 23112 6400 23164 6452
rect 22192 6332 22244 6384
rect 22652 6332 22704 6384
rect 23572 6400 23624 6452
rect 25504 6443 25556 6452
rect 25504 6409 25513 6443
rect 25513 6409 25547 6443
rect 25547 6409 25556 6443
rect 25504 6400 25556 6409
rect 25780 6400 25832 6452
rect 26332 6400 26384 6452
rect 27620 6400 27672 6452
rect 28816 6400 28868 6452
rect 29092 6400 29144 6452
rect 24308 6332 24360 6384
rect 25320 6332 25372 6384
rect 20720 6196 20772 6248
rect 20812 6196 20864 6248
rect 22192 6239 22244 6248
rect 22192 6205 22201 6239
rect 22201 6205 22235 6239
rect 22235 6205 22244 6239
rect 22192 6196 22244 6205
rect 26608 6264 26660 6316
rect 27896 6332 27948 6384
rect 27436 6264 27488 6316
rect 25780 6128 25832 6180
rect 28540 6196 28592 6248
rect 29092 6196 29144 6248
rect 27160 6128 27212 6180
rect 27712 6128 27764 6180
rect 23572 6060 23624 6112
rect 26240 6103 26292 6112
rect 26240 6069 26249 6103
rect 26249 6069 26283 6103
rect 26283 6069 26292 6103
rect 26240 6060 26292 6069
rect 26516 6103 26568 6112
rect 26516 6069 26525 6103
rect 26525 6069 26559 6103
rect 26559 6069 26568 6103
rect 26516 6060 26568 6069
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 23480 5856 23532 5908
rect 23572 5856 23624 5908
rect 23664 5763 23716 5772
rect 23664 5729 23673 5763
rect 23673 5729 23707 5763
rect 23707 5729 23716 5763
rect 23664 5720 23716 5729
rect 25688 5856 25740 5908
rect 26608 5856 26660 5908
rect 27988 5899 28040 5908
rect 27988 5865 27997 5899
rect 27997 5865 28031 5899
rect 28031 5865 28040 5899
rect 27988 5856 28040 5865
rect 28448 5856 28500 5908
rect 29092 5856 29144 5908
rect 27068 5720 27120 5772
rect 22652 5652 22704 5704
rect 25780 5652 25832 5704
rect 27896 5652 27948 5704
rect 28816 5695 28868 5704
rect 28816 5661 28825 5695
rect 28825 5661 28859 5695
rect 28859 5661 28868 5695
rect 28816 5652 28868 5661
rect 26516 5627 26568 5636
rect 26516 5593 26525 5627
rect 26525 5593 26559 5627
rect 26559 5593 26568 5627
rect 26516 5584 26568 5593
rect 26700 5516 26752 5568
rect 28172 5559 28224 5568
rect 28172 5525 28181 5559
rect 28181 5525 28215 5559
rect 28215 5525 28224 5559
rect 28172 5516 28224 5525
rect 29092 5559 29144 5568
rect 29092 5525 29101 5559
rect 29101 5525 29135 5559
rect 29135 5525 29144 5559
rect 29092 5516 29144 5525
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 35594 5414 35646 5466
rect 35658 5414 35710 5466
rect 35722 5414 35774 5466
rect 35786 5414 35838 5466
rect 35850 5414 35902 5466
rect 22192 5312 22244 5364
rect 24400 5312 24452 5364
rect 26240 5312 26292 5364
rect 26516 5312 26568 5364
rect 28172 5312 28224 5364
rect 29092 5312 29144 5364
rect 27988 5176 28040 5228
rect 26424 5151 26476 5160
rect 26424 5117 26433 5151
rect 26433 5117 26467 5151
rect 26467 5117 26476 5151
rect 26424 5108 26476 5117
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 26424 4768 26476 4820
rect 28356 4768 28408 4820
rect 27160 4564 27212 4616
rect 27436 4607 27488 4616
rect 27436 4573 27445 4607
rect 27445 4573 27479 4607
rect 27479 4573 27488 4607
rect 27436 4564 27488 4573
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 35594 4326 35646 4378
rect 35658 4326 35710 4378
rect 35722 4326 35774 4378
rect 35786 4326 35838 4378
rect 35850 4326 35902 4378
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 35594 3238 35646 3290
rect 35658 3238 35710 3290
rect 35722 3238 35774 3290
rect 35786 3238 35838 3290
rect 35850 3238 35902 3290
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 24216 2592 24268 2644
rect 23848 2388 23900 2440
rect 20 2320 72 2372
rect 11796 2363 11848 2372
rect 11796 2329 11805 2363
rect 11805 2329 11839 2363
rect 11839 2329 11848 2363
rect 11796 2320 11848 2329
rect 22100 2320 22152 2372
rect 18696 2252 18748 2304
rect 22008 2252 22060 2304
rect 35440 2252 35492 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 35594 2150 35646 2202
rect 35658 2150 35710 2202
rect 35722 2150 35774 2202
rect 35786 2150 35838 2202
rect 35850 2150 35902 2202
<< metal2 >>
rect 9678 39200 9734 40000
rect 21914 39200 21970 40000
rect 33506 39200 33562 40000
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 938 37496 994 37505
rect 4214 37499 4522 37508
rect 9692 37466 9720 39200
rect 938 37431 940 37440
rect 992 37431 994 37440
rect 9680 37460 9732 37466
rect 940 37402 992 37408
rect 9680 37402 9732 37408
rect 21928 37330 21956 39200
rect 21916 37324 21968 37330
rect 21916 37266 21968 37272
rect 33520 37262 33548 39200
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 22284 37256 22336 37262
rect 22284 37198 22336 37204
rect 33508 37256 33560 37262
rect 33508 37198 33560 37204
rect 10140 37188 10192 37194
rect 10140 37130 10192 37136
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 938 25256 994 25265
rect 938 25191 940 25200
rect 992 25191 994 25200
rect 940 25162 992 25168
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 10152 13530 10180 37130
rect 22296 26234 22324 37198
rect 26240 37188 26292 37194
rect 26240 37130 26292 37136
rect 22204 26206 22324 26234
rect 19616 25152 19668 25158
rect 19616 25094 19668 25100
rect 18972 15020 19024 15026
rect 18972 14962 19024 14968
rect 18788 14816 18840 14822
rect 18788 14758 18840 14764
rect 18800 14006 18828 14758
rect 18984 14618 19012 14962
rect 18972 14612 19024 14618
rect 18972 14554 19024 14560
rect 19628 14414 19656 25094
rect 22204 15586 22232 26206
rect 23664 16108 23716 16114
rect 23664 16050 23716 16056
rect 22376 16040 22428 16046
rect 22376 15982 22428 15988
rect 22284 15904 22336 15910
rect 22284 15846 22336 15852
rect 22296 15706 22324 15846
rect 22284 15700 22336 15706
rect 22284 15642 22336 15648
rect 22204 15570 22324 15586
rect 22204 15564 22336 15570
rect 22204 15558 22284 15564
rect 21088 15496 21140 15502
rect 21088 15438 21140 15444
rect 21916 15496 21968 15502
rect 21916 15438 21968 15444
rect 20536 15360 20588 15366
rect 20536 15302 20588 15308
rect 20548 15162 20576 15302
rect 21100 15162 21128 15438
rect 21180 15360 21232 15366
rect 21180 15302 21232 15308
rect 20536 15156 20588 15162
rect 20536 15098 20588 15104
rect 21088 15156 21140 15162
rect 21088 15098 21140 15104
rect 20536 14952 20588 14958
rect 20536 14894 20588 14900
rect 20548 14482 20576 14894
rect 20720 14816 20772 14822
rect 20720 14758 20772 14764
rect 20732 14618 20760 14758
rect 20720 14612 20772 14618
rect 20720 14554 20772 14560
rect 20076 14476 20128 14482
rect 20076 14418 20128 14424
rect 20536 14476 20588 14482
rect 20536 14418 20588 14424
rect 19616 14408 19668 14414
rect 19616 14350 19668 14356
rect 18788 14000 18840 14006
rect 18788 13942 18840 13948
rect 18604 13864 18656 13870
rect 18604 13806 18656 13812
rect 10140 13524 10192 13530
rect 10140 13466 10192 13472
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1412 12345 1440 12786
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 1398 12336 1454 12345
rect 18616 12306 18644 13806
rect 19628 13394 19656 14350
rect 19708 14272 19760 14278
rect 19708 14214 19760 14220
rect 19720 14074 19748 14214
rect 19708 14068 19760 14074
rect 19708 14010 19760 14016
rect 19616 13388 19668 13394
rect 19616 13330 19668 13336
rect 19432 13320 19484 13326
rect 19432 13262 19484 13268
rect 1398 12271 1454 12280
rect 18604 12300 18656 12306
rect 18604 12242 18656 12248
rect 18236 12096 18288 12102
rect 18236 12038 18288 12044
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 18248 11898 18276 12038
rect 18616 11898 18644 12242
rect 19444 12170 19472 13262
rect 19984 13184 20036 13190
rect 19984 13126 20036 13132
rect 19996 12918 20024 13126
rect 19984 12912 20036 12918
rect 19984 12854 20036 12860
rect 20088 12782 20116 14418
rect 20628 14000 20680 14006
rect 20628 13942 20680 13948
rect 20076 12776 20128 12782
rect 20076 12718 20128 12724
rect 19524 12640 19576 12646
rect 19524 12582 19576 12588
rect 19536 12170 19564 12582
rect 19984 12436 20036 12442
rect 20088 12434 20116 12718
rect 20036 12406 20116 12434
rect 19984 12378 20036 12384
rect 20640 12238 20668 13942
rect 20732 13326 20760 14554
rect 21192 14346 21220 15302
rect 21928 14958 21956 15438
rect 22204 15162 22232 15558
rect 22284 15506 22336 15512
rect 22192 15156 22244 15162
rect 22192 15098 22244 15104
rect 22284 15020 22336 15026
rect 22284 14962 22336 14968
rect 21916 14952 21968 14958
rect 21916 14894 21968 14900
rect 21916 14476 21968 14482
rect 21916 14418 21968 14424
rect 21180 14340 21232 14346
rect 21180 14282 21232 14288
rect 21928 14006 21956 14418
rect 22192 14408 22244 14414
rect 22112 14368 22192 14396
rect 21916 14000 21968 14006
rect 21916 13942 21968 13948
rect 20904 13932 20956 13938
rect 20904 13874 20956 13880
rect 20916 13462 20944 13874
rect 21916 13864 21968 13870
rect 21916 13806 21968 13812
rect 21928 13530 21956 13806
rect 21916 13524 21968 13530
rect 21916 13466 21968 13472
rect 20904 13456 20956 13462
rect 20904 13398 20956 13404
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 20732 12434 20760 13262
rect 21180 13252 21232 13258
rect 21180 13194 21232 13200
rect 21192 12986 21220 13194
rect 22008 13184 22060 13190
rect 22008 13126 22060 13132
rect 21180 12980 21232 12986
rect 21180 12922 21232 12928
rect 21456 12844 21508 12850
rect 21456 12786 21508 12792
rect 21088 12776 21140 12782
rect 21088 12718 21140 12724
rect 21100 12442 21128 12718
rect 21468 12442 21496 12786
rect 21088 12436 21140 12442
rect 20732 12406 20852 12434
rect 20824 12306 20852 12406
rect 21088 12378 21140 12384
rect 21456 12436 21508 12442
rect 21456 12378 21508 12384
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 20628 12232 20680 12238
rect 20628 12174 20680 12180
rect 19432 12164 19484 12170
rect 19432 12106 19484 12112
rect 19524 12164 19576 12170
rect 19524 12106 19576 12112
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18788 12096 18840 12102
rect 18788 12038 18840 12044
rect 18236 11892 18288 11898
rect 18236 11834 18288 11840
rect 18604 11892 18656 11898
rect 18604 11834 18656 11840
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 20 2372 72 2378
rect 20 2314 72 2320
rect 11796 2372 11848 2378
rect 11796 2314 11848 2320
rect 32 800 60 2314
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 11808 1170 11836 2314
rect 18708 2310 18736 12038
rect 18800 11354 18828 12038
rect 20442 11928 20498 11937
rect 20442 11863 20444 11872
rect 20496 11863 20498 11872
rect 20444 11834 20496 11840
rect 18788 11348 18840 11354
rect 18788 11290 18840 11296
rect 20456 11218 20484 11834
rect 20640 11830 20668 12174
rect 20628 11824 20680 11830
rect 20628 11766 20680 11772
rect 20444 11212 20496 11218
rect 20444 11154 20496 11160
rect 20640 11150 20668 11766
rect 20824 11626 20852 12242
rect 22020 12238 22048 13126
rect 22008 12232 22060 12238
rect 22008 12174 22060 12180
rect 20812 11620 20864 11626
rect 20812 11562 20864 11568
rect 20824 11354 20852 11562
rect 21824 11552 21876 11558
rect 21824 11494 21876 11500
rect 20812 11348 20864 11354
rect 20812 11290 20864 11296
rect 20628 11144 20680 11150
rect 20628 11086 20680 11092
rect 20824 10674 20852 11290
rect 20996 11076 21048 11082
rect 20996 11018 21048 11024
rect 21008 10810 21036 11018
rect 21836 10810 21864 11494
rect 20996 10804 21048 10810
rect 20996 10746 21048 10752
rect 21824 10804 21876 10810
rect 21824 10746 21876 10752
rect 20812 10668 20864 10674
rect 20812 10610 20864 10616
rect 20824 10266 20852 10610
rect 20812 10260 20864 10266
rect 20812 10202 20864 10208
rect 21732 9376 21784 9382
rect 21732 9318 21784 9324
rect 21456 8900 21508 8906
rect 21456 8842 21508 8848
rect 21468 8634 21496 8842
rect 21744 8634 21772 9318
rect 21824 9036 21876 9042
rect 21824 8978 21876 8984
rect 21456 8628 21508 8634
rect 21456 8570 21508 8576
rect 21732 8628 21784 8634
rect 21732 8570 21784 8576
rect 21836 8498 21864 8978
rect 21824 8492 21876 8498
rect 21824 8434 21876 8440
rect 21836 8090 21864 8434
rect 20812 8084 20864 8090
rect 20812 8026 20864 8032
rect 21824 8084 21876 8090
rect 21824 8026 21876 8032
rect 20536 7200 20588 7206
rect 20536 7142 20588 7148
rect 20548 7002 20576 7142
rect 20536 6996 20588 7002
rect 20536 6938 20588 6944
rect 20824 6866 20852 8026
rect 21824 7200 21876 7206
rect 21824 7142 21876 7148
rect 20812 6860 20864 6866
rect 20812 6802 20864 6808
rect 20720 6656 20772 6662
rect 20720 6598 20772 6604
rect 20732 6254 20760 6598
rect 20824 6458 20852 6802
rect 21836 6662 21864 7142
rect 21824 6656 21876 6662
rect 21824 6598 21876 6604
rect 20812 6452 20864 6458
rect 20812 6394 20864 6400
rect 20824 6254 20852 6394
rect 20720 6248 20772 6254
rect 20720 6190 20772 6196
rect 20812 6248 20864 6254
rect 20812 6190 20864 6196
rect 22020 2310 22048 12174
rect 22112 11830 22140 14368
rect 22192 14350 22244 14356
rect 22296 14278 22324 14962
rect 22388 14618 22416 15982
rect 22928 15496 22980 15502
rect 22928 15438 22980 15444
rect 22468 15360 22520 15366
rect 22468 15302 22520 15308
rect 22480 15162 22508 15302
rect 22468 15156 22520 15162
rect 22468 15098 22520 15104
rect 22940 14958 22968 15438
rect 23676 15162 23704 16050
rect 24216 16040 24268 16046
rect 24216 15982 24268 15988
rect 23940 15904 23992 15910
rect 23940 15846 23992 15852
rect 23952 15706 23980 15846
rect 23940 15700 23992 15706
rect 23940 15642 23992 15648
rect 23664 15156 23716 15162
rect 23664 15098 23716 15104
rect 22928 14952 22980 14958
rect 22928 14894 22980 14900
rect 24032 14952 24084 14958
rect 24032 14894 24084 14900
rect 22836 14816 22888 14822
rect 22836 14758 22888 14764
rect 22376 14612 22428 14618
rect 22376 14554 22428 14560
rect 22284 14272 22336 14278
rect 22284 14214 22336 14220
rect 22296 14074 22324 14214
rect 22284 14068 22336 14074
rect 22284 14010 22336 14016
rect 22192 13728 22244 13734
rect 22192 13670 22244 13676
rect 22204 12986 22232 13670
rect 22296 13326 22324 14010
rect 22284 13320 22336 13326
rect 22284 13262 22336 13268
rect 22192 12980 22244 12986
rect 22192 12922 22244 12928
rect 22388 12782 22416 14554
rect 22848 14482 22876 14758
rect 22836 14476 22888 14482
rect 22836 14418 22888 14424
rect 22940 14362 22968 14894
rect 24044 14482 24072 14894
rect 24032 14476 24084 14482
rect 24032 14418 24084 14424
rect 22848 14334 22968 14362
rect 22848 12850 22876 14334
rect 23664 14272 23716 14278
rect 23664 14214 23716 14220
rect 23676 14006 23704 14214
rect 23664 14000 23716 14006
rect 23584 13960 23664 13988
rect 23204 13864 23256 13870
rect 23204 13806 23256 13812
rect 23216 13530 23244 13806
rect 23204 13524 23256 13530
rect 23204 13466 23256 13472
rect 22928 13184 22980 13190
rect 22928 13126 22980 13132
rect 22836 12844 22888 12850
rect 22836 12786 22888 12792
rect 22376 12776 22428 12782
rect 22376 12718 22428 12724
rect 22560 12708 22612 12714
rect 22560 12650 22612 12656
rect 22100 11824 22152 11830
rect 22100 11766 22152 11772
rect 22112 11354 22140 11766
rect 22192 11756 22244 11762
rect 22192 11698 22244 11704
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 22204 11218 22232 11698
rect 22572 11694 22600 12650
rect 22940 12646 22968 13126
rect 23204 12776 23256 12782
rect 23204 12718 23256 12724
rect 22928 12640 22980 12646
rect 22928 12582 22980 12588
rect 22940 12306 22968 12582
rect 22928 12300 22980 12306
rect 22928 12242 22980 12248
rect 23216 11830 23244 12718
rect 23584 11830 23612 13960
rect 23664 13942 23716 13948
rect 24044 13530 24072 14418
rect 24032 13524 24084 13530
rect 24032 13466 24084 13472
rect 24044 13394 24072 13466
rect 24228 13394 24256 15982
rect 24952 15360 25004 15366
rect 24952 15302 25004 15308
rect 24964 15162 24992 15302
rect 24952 15156 25004 15162
rect 24952 15098 25004 15104
rect 24492 15020 24544 15026
rect 24492 14962 24544 14968
rect 25412 15020 25464 15026
rect 25412 14962 25464 14968
rect 24400 14272 24452 14278
rect 24400 14214 24452 14220
rect 24412 13394 24440 14214
rect 24504 13870 24532 14962
rect 25044 14816 25096 14822
rect 25044 14758 25096 14764
rect 25320 14816 25372 14822
rect 25320 14758 25372 14764
rect 25056 14550 25084 14758
rect 25044 14544 25096 14550
rect 25044 14486 25096 14492
rect 24492 13864 24544 13870
rect 24492 13806 24544 13812
rect 24860 13864 24912 13870
rect 24860 13806 24912 13812
rect 24872 13394 24900 13806
rect 24032 13388 24084 13394
rect 24032 13330 24084 13336
rect 24216 13388 24268 13394
rect 24216 13330 24268 13336
rect 24400 13388 24452 13394
rect 24400 13330 24452 13336
rect 24860 13388 24912 13394
rect 24860 13330 24912 13336
rect 23664 12640 23716 12646
rect 23664 12582 23716 12588
rect 23756 12640 23808 12646
rect 23756 12582 23808 12588
rect 23676 12442 23704 12582
rect 23664 12436 23716 12442
rect 23768 12434 23796 12582
rect 23768 12406 23888 12434
rect 23664 12378 23716 12384
rect 23860 12238 23888 12406
rect 23848 12232 23900 12238
rect 23848 12174 23900 12180
rect 23204 11824 23256 11830
rect 23572 11824 23624 11830
rect 23204 11766 23256 11772
rect 23400 11784 23572 11812
rect 22560 11688 22612 11694
rect 22560 11630 22612 11636
rect 22928 11688 22980 11694
rect 22928 11630 22980 11636
rect 22192 11212 22244 11218
rect 22192 11154 22244 11160
rect 22940 11082 22968 11630
rect 23112 11552 23164 11558
rect 23112 11494 23164 11500
rect 23020 11348 23072 11354
rect 23020 11290 23072 11296
rect 22928 11076 22980 11082
rect 22928 11018 22980 11024
rect 22836 11008 22888 11014
rect 22836 10950 22888 10956
rect 22848 10810 22876 10950
rect 22836 10804 22888 10810
rect 22836 10746 22888 10752
rect 22468 10464 22520 10470
rect 22468 10406 22520 10412
rect 22480 9994 22508 10406
rect 22940 9994 22968 11018
rect 22468 9988 22520 9994
rect 22468 9930 22520 9936
rect 22928 9988 22980 9994
rect 22928 9930 22980 9936
rect 22100 8424 22152 8430
rect 22100 8366 22152 8372
rect 22112 8090 22140 8366
rect 22100 8084 22152 8090
rect 22100 8026 22152 8032
rect 22480 7886 22508 9930
rect 22744 9920 22796 9926
rect 22744 9862 22796 9868
rect 22756 9586 22784 9862
rect 23032 9654 23060 11290
rect 23124 11098 23152 11494
rect 23216 11286 23244 11766
rect 23204 11280 23256 11286
rect 23204 11222 23256 11228
rect 23124 11082 23244 11098
rect 23124 11076 23256 11082
rect 23124 11070 23204 11076
rect 23204 11018 23256 11024
rect 23400 10742 23428 11784
rect 23572 11766 23624 11772
rect 23756 11688 23808 11694
rect 23756 11630 23808 11636
rect 23572 11280 23624 11286
rect 23572 11222 23624 11228
rect 23480 11008 23532 11014
rect 23480 10950 23532 10956
rect 23388 10736 23440 10742
rect 23388 10678 23440 10684
rect 23492 10266 23520 10950
rect 23584 10810 23612 11222
rect 23768 10810 23796 11630
rect 23848 11144 23900 11150
rect 23848 11086 23900 11092
rect 23860 10810 23888 11086
rect 23940 11008 23992 11014
rect 23940 10950 23992 10956
rect 23572 10804 23624 10810
rect 23572 10746 23624 10752
rect 23756 10804 23808 10810
rect 23756 10746 23808 10752
rect 23848 10804 23900 10810
rect 23848 10746 23900 10752
rect 23952 10674 23980 10950
rect 23940 10668 23992 10674
rect 23940 10610 23992 10616
rect 23480 10260 23532 10266
rect 23480 10202 23532 10208
rect 23296 10056 23348 10062
rect 23296 9998 23348 10004
rect 23020 9648 23072 9654
rect 23020 9590 23072 9596
rect 22744 9580 22796 9586
rect 22744 9522 22796 9528
rect 22836 9376 22888 9382
rect 22836 9318 22888 9324
rect 22848 9042 22876 9318
rect 23032 9194 23060 9590
rect 22940 9166 23060 9194
rect 23308 9178 23336 9998
rect 23296 9172 23348 9178
rect 22836 9036 22888 9042
rect 22836 8978 22888 8984
rect 22940 8974 22968 9166
rect 23296 9114 23348 9120
rect 23020 9036 23072 9042
rect 23020 8978 23072 8984
rect 22560 8968 22612 8974
rect 22560 8910 22612 8916
rect 22928 8968 22980 8974
rect 22928 8910 22980 8916
rect 22572 8566 22600 8910
rect 22560 8560 22612 8566
rect 22560 8502 22612 8508
rect 22468 7880 22520 7886
rect 22468 7822 22520 7828
rect 22572 6798 22600 8502
rect 23032 7886 23060 8978
rect 23308 8090 23336 9114
rect 24032 8424 24084 8430
rect 24032 8366 24084 8372
rect 23572 8288 23624 8294
rect 23572 8230 23624 8236
rect 23664 8288 23716 8294
rect 23664 8230 23716 8236
rect 23296 8084 23348 8090
rect 23296 8026 23348 8032
rect 23584 7954 23612 8230
rect 23676 8090 23704 8230
rect 24044 8090 24072 8366
rect 23664 8084 23716 8090
rect 23664 8026 23716 8032
rect 24032 8084 24084 8090
rect 24032 8026 24084 8032
rect 23572 7948 23624 7954
rect 23572 7890 23624 7896
rect 23020 7880 23072 7886
rect 23020 7822 23072 7828
rect 22928 7812 22980 7818
rect 22928 7754 22980 7760
rect 22940 7546 22968 7754
rect 22928 7540 22980 7546
rect 22928 7482 22980 7488
rect 23848 7404 23900 7410
rect 23848 7346 23900 7352
rect 22744 7336 22796 7342
rect 22744 7278 22796 7284
rect 23020 7336 23072 7342
rect 23020 7278 23072 7284
rect 23664 7336 23716 7342
rect 23664 7278 23716 7284
rect 22756 6866 22784 7278
rect 22744 6860 22796 6866
rect 22744 6802 22796 6808
rect 22192 6792 22244 6798
rect 22192 6734 22244 6740
rect 22560 6792 22612 6798
rect 22560 6734 22612 6740
rect 22100 6724 22152 6730
rect 22100 6666 22152 6672
rect 22112 2378 22140 6666
rect 22204 6390 22232 6734
rect 23032 6458 23060 7278
rect 23676 6866 23704 7278
rect 23860 6866 23888 7346
rect 24124 7200 24176 7206
rect 24124 7142 24176 7148
rect 23480 6860 23532 6866
rect 23480 6802 23532 6808
rect 23664 6860 23716 6866
rect 23664 6802 23716 6808
rect 23848 6860 23900 6866
rect 23848 6802 23900 6808
rect 23112 6724 23164 6730
rect 23112 6666 23164 6672
rect 23124 6458 23152 6666
rect 23020 6452 23072 6458
rect 23020 6394 23072 6400
rect 23112 6452 23164 6458
rect 23112 6394 23164 6400
rect 22192 6384 22244 6390
rect 22192 6326 22244 6332
rect 22652 6384 22704 6390
rect 22652 6326 22704 6332
rect 22192 6248 22244 6254
rect 22192 6190 22244 6196
rect 22204 5370 22232 6190
rect 22664 5710 22692 6326
rect 23492 5914 23520 6802
rect 23676 6746 23704 6802
rect 24136 6798 24164 7142
rect 23584 6718 23704 6746
rect 24124 6792 24176 6798
rect 24124 6734 24176 6740
rect 23584 6458 23612 6718
rect 23664 6656 23716 6662
rect 23664 6598 23716 6604
rect 23572 6452 23624 6458
rect 23572 6394 23624 6400
rect 23572 6112 23624 6118
rect 23572 6054 23624 6060
rect 23584 5914 23612 6054
rect 23480 5908 23532 5914
rect 23480 5850 23532 5856
rect 23572 5908 23624 5914
rect 23572 5850 23624 5856
rect 23676 5778 23704 6598
rect 23664 5772 23716 5778
rect 23664 5714 23716 5720
rect 22652 5704 22704 5710
rect 22652 5646 22704 5652
rect 22192 5364 22244 5370
rect 22192 5306 22244 5312
rect 24228 2650 24256 13330
rect 24400 12844 24452 12850
rect 24400 12786 24452 12792
rect 24412 12646 24440 12786
rect 25056 12782 25084 14486
rect 25332 14414 25360 14758
rect 25228 14408 25280 14414
rect 25228 14350 25280 14356
rect 25320 14408 25372 14414
rect 25320 14350 25372 14356
rect 25240 13734 25268 14350
rect 25424 14346 25452 14962
rect 25504 14816 25556 14822
rect 25504 14758 25556 14764
rect 25412 14340 25464 14346
rect 25412 14282 25464 14288
rect 25516 14074 25544 14758
rect 26252 14482 26280 37130
rect 33692 37120 33744 37126
rect 33692 37062 33744 37068
rect 33704 16114 33732 37062
rect 35594 37020 35902 37029
rect 35594 37018 35600 37020
rect 35656 37018 35680 37020
rect 35736 37018 35760 37020
rect 35816 37018 35840 37020
rect 35896 37018 35902 37020
rect 35656 36966 35658 37018
rect 35838 36966 35840 37018
rect 35594 36964 35600 36966
rect 35656 36964 35680 36966
rect 35736 36964 35760 36966
rect 35816 36964 35840 36966
rect 35896 36964 35902 36966
rect 35594 36955 35902 36964
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 35594 35932 35902 35941
rect 35594 35930 35600 35932
rect 35656 35930 35680 35932
rect 35736 35930 35760 35932
rect 35816 35930 35840 35932
rect 35896 35930 35902 35932
rect 35656 35878 35658 35930
rect 35838 35878 35840 35930
rect 35594 35876 35600 35878
rect 35656 35876 35680 35878
rect 35736 35876 35760 35878
rect 35816 35876 35840 35878
rect 35896 35876 35902 35878
rect 35594 35867 35902 35876
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 35594 34844 35902 34853
rect 35594 34842 35600 34844
rect 35656 34842 35680 34844
rect 35736 34842 35760 34844
rect 35816 34842 35840 34844
rect 35896 34842 35902 34844
rect 35656 34790 35658 34842
rect 35838 34790 35840 34842
rect 35594 34788 35600 34790
rect 35656 34788 35680 34790
rect 35736 34788 35760 34790
rect 35816 34788 35840 34790
rect 35896 34788 35902 34790
rect 35594 34779 35902 34788
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 35594 33756 35902 33765
rect 35594 33754 35600 33756
rect 35656 33754 35680 33756
rect 35736 33754 35760 33756
rect 35816 33754 35840 33756
rect 35896 33754 35902 33756
rect 35656 33702 35658 33754
rect 35838 33702 35840 33754
rect 35594 33700 35600 33702
rect 35656 33700 35680 33702
rect 35736 33700 35760 33702
rect 35816 33700 35840 33702
rect 35896 33700 35902 33702
rect 35594 33691 35902 33700
rect 38844 33516 38896 33522
rect 38844 33458 38896 33464
rect 38856 33425 38884 33458
rect 38842 33416 38898 33425
rect 38842 33351 38898 33360
rect 38292 33312 38344 33318
rect 38292 33254 38344 33260
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 35594 32668 35902 32677
rect 35594 32666 35600 32668
rect 35656 32666 35680 32668
rect 35736 32666 35760 32668
rect 35816 32666 35840 32668
rect 35896 32666 35902 32668
rect 35656 32614 35658 32666
rect 35838 32614 35840 32666
rect 35594 32612 35600 32614
rect 35656 32612 35680 32614
rect 35736 32612 35760 32614
rect 35816 32612 35840 32614
rect 35896 32612 35902 32614
rect 35594 32603 35902 32612
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 35594 31580 35902 31589
rect 35594 31578 35600 31580
rect 35656 31578 35680 31580
rect 35736 31578 35760 31580
rect 35816 31578 35840 31580
rect 35896 31578 35902 31580
rect 35656 31526 35658 31578
rect 35838 31526 35840 31578
rect 35594 31524 35600 31526
rect 35656 31524 35680 31526
rect 35736 31524 35760 31526
rect 35816 31524 35840 31526
rect 35896 31524 35902 31526
rect 35594 31515 35902 31524
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 35594 30492 35902 30501
rect 35594 30490 35600 30492
rect 35656 30490 35680 30492
rect 35736 30490 35760 30492
rect 35816 30490 35840 30492
rect 35896 30490 35902 30492
rect 35656 30438 35658 30490
rect 35838 30438 35840 30490
rect 35594 30436 35600 30438
rect 35656 30436 35680 30438
rect 35736 30436 35760 30438
rect 35816 30436 35840 30438
rect 35896 30436 35902 30438
rect 35594 30427 35902 30436
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 35594 29404 35902 29413
rect 35594 29402 35600 29404
rect 35656 29402 35680 29404
rect 35736 29402 35760 29404
rect 35816 29402 35840 29404
rect 35896 29402 35902 29404
rect 35656 29350 35658 29402
rect 35838 29350 35840 29402
rect 35594 29348 35600 29350
rect 35656 29348 35680 29350
rect 35736 29348 35760 29350
rect 35816 29348 35840 29350
rect 35896 29348 35902 29350
rect 35594 29339 35902 29348
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 35594 28316 35902 28325
rect 35594 28314 35600 28316
rect 35656 28314 35680 28316
rect 35736 28314 35760 28316
rect 35816 28314 35840 28316
rect 35896 28314 35902 28316
rect 35656 28262 35658 28314
rect 35838 28262 35840 28314
rect 35594 28260 35600 28262
rect 35656 28260 35680 28262
rect 35736 28260 35760 28262
rect 35816 28260 35840 28262
rect 35896 28260 35902 28262
rect 35594 28251 35902 28260
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35594 27228 35902 27237
rect 35594 27226 35600 27228
rect 35656 27226 35680 27228
rect 35736 27226 35760 27228
rect 35816 27226 35840 27228
rect 35896 27226 35902 27228
rect 35656 27174 35658 27226
rect 35838 27174 35840 27226
rect 35594 27172 35600 27174
rect 35656 27172 35680 27174
rect 35736 27172 35760 27174
rect 35816 27172 35840 27174
rect 35896 27172 35902 27174
rect 35594 27163 35902 27172
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35594 26140 35902 26149
rect 35594 26138 35600 26140
rect 35656 26138 35680 26140
rect 35736 26138 35760 26140
rect 35816 26138 35840 26140
rect 35896 26138 35902 26140
rect 35656 26086 35658 26138
rect 35838 26086 35840 26138
rect 35594 26084 35600 26086
rect 35656 26084 35680 26086
rect 35736 26084 35760 26086
rect 35816 26084 35840 26086
rect 35896 26084 35902 26086
rect 35594 26075 35902 26084
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 35594 25052 35902 25061
rect 35594 25050 35600 25052
rect 35656 25050 35680 25052
rect 35736 25050 35760 25052
rect 35816 25050 35840 25052
rect 35896 25050 35902 25052
rect 35656 24998 35658 25050
rect 35838 24998 35840 25050
rect 35594 24996 35600 24998
rect 35656 24996 35680 24998
rect 35736 24996 35760 24998
rect 35816 24996 35840 24998
rect 35896 24996 35902 24998
rect 35594 24987 35902 24996
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35594 23964 35902 23973
rect 35594 23962 35600 23964
rect 35656 23962 35680 23964
rect 35736 23962 35760 23964
rect 35816 23962 35840 23964
rect 35896 23962 35902 23964
rect 35656 23910 35658 23962
rect 35838 23910 35840 23962
rect 35594 23908 35600 23910
rect 35656 23908 35680 23910
rect 35736 23908 35760 23910
rect 35816 23908 35840 23910
rect 35896 23908 35902 23910
rect 35594 23899 35902 23908
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 35594 22876 35902 22885
rect 35594 22874 35600 22876
rect 35656 22874 35680 22876
rect 35736 22874 35760 22876
rect 35816 22874 35840 22876
rect 35896 22874 35902 22876
rect 35656 22822 35658 22874
rect 35838 22822 35840 22874
rect 35594 22820 35600 22822
rect 35656 22820 35680 22822
rect 35736 22820 35760 22822
rect 35816 22820 35840 22822
rect 35896 22820 35902 22822
rect 35594 22811 35902 22820
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 35594 21788 35902 21797
rect 35594 21786 35600 21788
rect 35656 21786 35680 21788
rect 35736 21786 35760 21788
rect 35816 21786 35840 21788
rect 35896 21786 35902 21788
rect 35656 21734 35658 21786
rect 35838 21734 35840 21786
rect 35594 21732 35600 21734
rect 35656 21732 35680 21734
rect 35736 21732 35760 21734
rect 35816 21732 35840 21734
rect 35896 21732 35902 21734
rect 35594 21723 35902 21732
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 35594 20700 35902 20709
rect 35594 20698 35600 20700
rect 35656 20698 35680 20700
rect 35736 20698 35760 20700
rect 35816 20698 35840 20700
rect 35896 20698 35902 20700
rect 35656 20646 35658 20698
rect 35838 20646 35840 20698
rect 35594 20644 35600 20646
rect 35656 20644 35680 20646
rect 35736 20644 35760 20646
rect 35816 20644 35840 20646
rect 35896 20644 35902 20646
rect 35594 20635 35902 20644
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35594 19612 35902 19621
rect 35594 19610 35600 19612
rect 35656 19610 35680 19612
rect 35736 19610 35760 19612
rect 35816 19610 35840 19612
rect 35896 19610 35902 19612
rect 35656 19558 35658 19610
rect 35838 19558 35840 19610
rect 35594 19556 35600 19558
rect 35656 19556 35680 19558
rect 35736 19556 35760 19558
rect 35816 19556 35840 19558
rect 35896 19556 35902 19558
rect 35594 19547 35902 19556
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 35594 18524 35902 18533
rect 35594 18522 35600 18524
rect 35656 18522 35680 18524
rect 35736 18522 35760 18524
rect 35816 18522 35840 18524
rect 35896 18522 35902 18524
rect 35656 18470 35658 18522
rect 35838 18470 35840 18522
rect 35594 18468 35600 18470
rect 35656 18468 35680 18470
rect 35736 18468 35760 18470
rect 35816 18468 35840 18470
rect 35896 18468 35902 18470
rect 35594 18459 35902 18468
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35594 17436 35902 17445
rect 35594 17434 35600 17436
rect 35656 17434 35680 17436
rect 35736 17434 35760 17436
rect 35816 17434 35840 17436
rect 35896 17434 35902 17436
rect 35656 17382 35658 17434
rect 35838 17382 35840 17434
rect 35594 17380 35600 17382
rect 35656 17380 35680 17382
rect 35736 17380 35760 17382
rect 35816 17380 35840 17382
rect 35896 17380 35902 17382
rect 35594 17371 35902 17380
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35594 16348 35902 16357
rect 35594 16346 35600 16348
rect 35656 16346 35680 16348
rect 35736 16346 35760 16348
rect 35816 16346 35840 16348
rect 35896 16346 35902 16348
rect 35656 16294 35658 16346
rect 35838 16294 35840 16346
rect 35594 16292 35600 16294
rect 35656 16292 35680 16294
rect 35736 16292 35760 16294
rect 35816 16292 35840 16294
rect 35896 16292 35902 16294
rect 35594 16283 35902 16292
rect 33692 16108 33744 16114
rect 33692 16050 33744 16056
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 38304 15502 38332 33254
rect 38292 15496 38344 15502
rect 38292 15438 38344 15444
rect 35594 15260 35902 15269
rect 35594 15258 35600 15260
rect 35656 15258 35680 15260
rect 35736 15258 35760 15260
rect 35816 15258 35840 15260
rect 35896 15258 35902 15260
rect 35656 15206 35658 15258
rect 35838 15206 35840 15258
rect 35594 15204 35600 15206
rect 35656 15204 35680 15206
rect 35736 15204 35760 15206
rect 35816 15204 35840 15206
rect 35896 15204 35902 15206
rect 35594 15195 35902 15204
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 26240 14476 26292 14482
rect 26240 14418 26292 14424
rect 27160 14476 27212 14482
rect 27160 14418 27212 14424
rect 27528 14476 27580 14482
rect 27528 14418 27580 14424
rect 25780 14272 25832 14278
rect 25780 14214 25832 14220
rect 25792 14074 25820 14214
rect 25504 14068 25556 14074
rect 25504 14010 25556 14016
rect 25780 14068 25832 14074
rect 25780 14010 25832 14016
rect 26700 14000 26752 14006
rect 26700 13942 26752 13948
rect 25872 13864 25924 13870
rect 25872 13806 25924 13812
rect 25228 13728 25280 13734
rect 25228 13670 25280 13676
rect 25240 12850 25268 13670
rect 25320 13320 25372 13326
rect 25320 13262 25372 13268
rect 25228 12844 25280 12850
rect 25228 12786 25280 12792
rect 24676 12776 24728 12782
rect 24676 12718 24728 12724
rect 25044 12776 25096 12782
rect 25044 12718 25096 12724
rect 24400 12640 24452 12646
rect 24400 12582 24452 12588
rect 24492 12640 24544 12646
rect 24492 12582 24544 12588
rect 24400 11144 24452 11150
rect 24400 11086 24452 11092
rect 24412 10130 24440 11086
rect 24504 10130 24532 12582
rect 24584 12096 24636 12102
rect 24584 12038 24636 12044
rect 24596 11558 24624 12038
rect 24688 11937 24716 12718
rect 24952 12708 25004 12714
rect 24952 12650 25004 12656
rect 24674 11928 24730 11937
rect 24674 11863 24730 11872
rect 24676 11824 24728 11830
rect 24676 11766 24728 11772
rect 24584 11552 24636 11558
rect 24584 11494 24636 11500
rect 24596 10130 24624 11494
rect 24688 11014 24716 11766
rect 24860 11552 24912 11558
rect 24860 11494 24912 11500
rect 24676 11008 24728 11014
rect 24676 10950 24728 10956
rect 24688 10538 24716 10950
rect 24872 10674 24900 11494
rect 24964 11150 24992 12650
rect 25228 12096 25280 12102
rect 25228 12038 25280 12044
rect 25136 11756 25188 11762
rect 25136 11698 25188 11704
rect 25044 11552 25096 11558
rect 25044 11494 25096 11500
rect 25056 11150 25084 11494
rect 25148 11218 25176 11698
rect 25240 11354 25268 12038
rect 25332 11354 25360 13262
rect 25504 12708 25556 12714
rect 25504 12650 25556 12656
rect 25412 12232 25464 12238
rect 25412 12174 25464 12180
rect 25228 11348 25280 11354
rect 25228 11290 25280 11296
rect 25320 11348 25372 11354
rect 25320 11290 25372 11296
rect 25424 11234 25452 12174
rect 25136 11212 25188 11218
rect 25136 11154 25188 11160
rect 25332 11206 25452 11234
rect 24952 11144 25004 11150
rect 24952 11086 25004 11092
rect 25044 11144 25096 11150
rect 25044 11086 25096 11092
rect 24860 10668 24912 10674
rect 24860 10610 24912 10616
rect 24676 10532 24728 10538
rect 24676 10474 24728 10480
rect 24964 10130 24992 11086
rect 24400 10124 24452 10130
rect 24400 10066 24452 10072
rect 24492 10124 24544 10130
rect 24492 10066 24544 10072
rect 24584 10124 24636 10130
rect 24584 10066 24636 10072
rect 24952 10124 25004 10130
rect 24952 10066 25004 10072
rect 24952 9920 25004 9926
rect 24952 9862 25004 9868
rect 24964 9722 24992 9862
rect 24952 9716 25004 9722
rect 24952 9658 25004 9664
rect 25056 9654 25084 11086
rect 25148 10266 25176 11154
rect 25332 11082 25360 11206
rect 25412 11144 25464 11150
rect 25410 11112 25412 11121
rect 25464 11112 25466 11121
rect 25320 11076 25372 11082
rect 25410 11047 25466 11056
rect 25320 11018 25372 11024
rect 25228 10804 25280 10810
rect 25228 10746 25280 10752
rect 25136 10260 25188 10266
rect 25136 10202 25188 10208
rect 25136 10124 25188 10130
rect 25136 10066 25188 10072
rect 24584 9648 24636 9654
rect 24504 9608 24584 9636
rect 24308 9512 24360 9518
rect 24308 9454 24360 9460
rect 24320 9178 24348 9454
rect 24308 9172 24360 9178
rect 24308 9114 24360 9120
rect 24504 8294 24532 9608
rect 24584 9590 24636 9596
rect 25044 9648 25096 9654
rect 25044 9590 25096 9596
rect 24676 9512 24728 9518
rect 24596 9460 24676 9466
rect 24596 9454 24728 9460
rect 24596 9438 24716 9454
rect 24596 9178 24624 9438
rect 24676 9376 24728 9382
rect 24676 9318 24728 9324
rect 24688 9178 24716 9318
rect 24584 9172 24636 9178
rect 24584 9114 24636 9120
rect 24676 9172 24728 9178
rect 24676 9114 24728 9120
rect 24492 8288 24544 8294
rect 24492 8230 24544 8236
rect 24504 7818 24532 8230
rect 24492 7812 24544 7818
rect 24492 7754 24544 7760
rect 24504 7478 24532 7754
rect 24492 7472 24544 7478
rect 24492 7414 24544 7420
rect 24400 7404 24452 7410
rect 24400 7346 24452 7352
rect 24308 7200 24360 7206
rect 24308 7142 24360 7148
rect 24320 6390 24348 7142
rect 24412 6798 24440 7346
rect 24504 6798 24532 7414
rect 24860 7404 24912 7410
rect 24860 7346 24912 7352
rect 24872 7002 24900 7346
rect 24860 6996 24912 7002
rect 24860 6938 24912 6944
rect 24400 6792 24452 6798
rect 24400 6734 24452 6740
rect 24492 6792 24544 6798
rect 24492 6734 24544 6740
rect 24400 6656 24452 6662
rect 24400 6598 24452 6604
rect 24308 6384 24360 6390
rect 24308 6326 24360 6332
rect 24412 5370 24440 6598
rect 25148 6474 25176 10066
rect 25240 9382 25268 10746
rect 25332 9382 25360 11018
rect 25424 10146 25452 11047
rect 25516 10266 25544 12650
rect 25884 12306 25912 13806
rect 26240 13252 26292 13258
rect 26240 13194 26292 13200
rect 26252 12986 26280 13194
rect 26608 13184 26660 13190
rect 26608 13126 26660 13132
rect 26240 12980 26292 12986
rect 26240 12922 26292 12928
rect 26252 12782 26280 12922
rect 25964 12776 26016 12782
rect 25964 12718 26016 12724
rect 26240 12776 26292 12782
rect 26240 12718 26292 12724
rect 26424 12776 26476 12782
rect 26424 12718 26476 12724
rect 25872 12300 25924 12306
rect 25872 12242 25924 12248
rect 25976 12238 26004 12718
rect 26332 12708 26384 12714
rect 26332 12650 26384 12656
rect 25964 12232 26016 12238
rect 25964 12174 26016 12180
rect 26240 12232 26292 12238
rect 26240 12174 26292 12180
rect 25964 12096 26016 12102
rect 25964 12038 26016 12044
rect 25596 11620 25648 11626
rect 25596 11562 25648 11568
rect 25608 11082 25636 11562
rect 25976 11354 26004 12038
rect 25964 11348 26016 11354
rect 25964 11290 26016 11296
rect 26148 11348 26200 11354
rect 26148 11290 26200 11296
rect 25596 11076 25648 11082
rect 25596 11018 25648 11024
rect 25872 11076 25924 11082
rect 25872 11018 25924 11024
rect 25884 10674 25912 11018
rect 25872 10668 25924 10674
rect 25872 10610 25924 10616
rect 25688 10600 25740 10606
rect 25688 10542 25740 10548
rect 25504 10260 25556 10266
rect 25504 10202 25556 10208
rect 25424 10118 25544 10146
rect 25412 10056 25464 10062
rect 25412 9998 25464 10004
rect 25424 9382 25452 9998
rect 25516 9926 25544 10118
rect 25504 9920 25556 9926
rect 25504 9862 25556 9868
rect 25596 9920 25648 9926
rect 25596 9862 25648 9868
rect 25516 9654 25544 9862
rect 25504 9648 25556 9654
rect 25504 9590 25556 9596
rect 25504 9444 25556 9450
rect 25504 9386 25556 9392
rect 25228 9376 25280 9382
rect 25228 9318 25280 9324
rect 25320 9376 25372 9382
rect 25320 9318 25372 9324
rect 25412 9376 25464 9382
rect 25412 9318 25464 9324
rect 25424 7750 25452 9318
rect 25516 9042 25544 9386
rect 25504 9036 25556 9042
rect 25504 8978 25556 8984
rect 25608 8838 25636 9862
rect 25700 9722 25728 10542
rect 25780 10056 25832 10062
rect 25780 9998 25832 10004
rect 25688 9716 25740 9722
rect 25688 9658 25740 9664
rect 25792 9602 25820 9998
rect 25884 9722 25912 10610
rect 25964 10464 26016 10470
rect 25964 10406 26016 10412
rect 25976 10062 26004 10406
rect 25964 10056 26016 10062
rect 26016 10004 26096 10010
rect 25964 9998 26096 10004
rect 25976 9982 26096 9998
rect 25964 9920 26016 9926
rect 25964 9862 26016 9868
rect 25872 9716 25924 9722
rect 25872 9658 25924 9664
rect 25976 9625 26004 9862
rect 25962 9616 26018 9625
rect 25792 9586 25912 9602
rect 25792 9580 25924 9586
rect 25792 9574 25872 9580
rect 25962 9551 26018 9560
rect 25872 9522 25924 9528
rect 25780 9172 25832 9178
rect 25780 9114 25832 9120
rect 25792 8906 25820 9114
rect 25780 8900 25832 8906
rect 25780 8842 25832 8848
rect 25596 8832 25648 8838
rect 25596 8774 25648 8780
rect 25792 8566 25820 8842
rect 25780 8560 25832 8566
rect 25780 8502 25832 8508
rect 25412 7744 25464 7750
rect 25412 7686 25464 7692
rect 25504 6792 25556 6798
rect 25504 6734 25556 6740
rect 25148 6446 25360 6474
rect 25516 6458 25544 6734
rect 25688 6656 25740 6662
rect 25688 6598 25740 6604
rect 25332 6390 25360 6446
rect 25504 6452 25556 6458
rect 25504 6394 25556 6400
rect 25320 6384 25372 6390
rect 25320 6326 25372 6332
rect 25700 5914 25728 6598
rect 25792 6458 25820 8502
rect 25884 7546 25912 9522
rect 25976 9518 26004 9551
rect 25964 9512 26016 9518
rect 25964 9454 26016 9460
rect 26068 7886 26096 9982
rect 26160 9722 26188 11290
rect 26252 11121 26280 12174
rect 26344 11762 26372 12650
rect 26436 12374 26464 12718
rect 26424 12368 26476 12374
rect 26424 12310 26476 12316
rect 26620 12306 26648 13126
rect 26608 12300 26660 12306
rect 26608 12242 26660 12248
rect 26424 12164 26476 12170
rect 26424 12106 26476 12112
rect 26436 11898 26464 12106
rect 26424 11892 26476 11898
rect 26424 11834 26476 11840
rect 26332 11756 26384 11762
rect 26332 11698 26384 11704
rect 26238 11112 26294 11121
rect 26238 11047 26294 11056
rect 26238 10976 26294 10985
rect 26238 10911 26294 10920
rect 26252 10742 26280 10911
rect 26344 10810 26372 11698
rect 26436 11642 26464 11834
rect 26436 11614 26556 11642
rect 26424 11552 26476 11558
rect 26424 11494 26476 11500
rect 26436 11014 26464 11494
rect 26528 11218 26556 11614
rect 26608 11552 26660 11558
rect 26608 11494 26660 11500
rect 26620 11286 26648 11494
rect 26608 11280 26660 11286
rect 26608 11222 26660 11228
rect 26516 11212 26568 11218
rect 26516 11154 26568 11160
rect 26712 11098 26740 13942
rect 27172 13258 27200 14418
rect 27344 14340 27396 14346
rect 27344 14282 27396 14288
rect 27160 13252 27212 13258
rect 27160 13194 27212 13200
rect 27356 12986 27384 14282
rect 27540 13326 27568 14418
rect 27896 14340 27948 14346
rect 27896 14282 27948 14288
rect 27908 14074 27936 14282
rect 35594 14172 35902 14181
rect 35594 14170 35600 14172
rect 35656 14170 35680 14172
rect 35736 14170 35760 14172
rect 35816 14170 35840 14172
rect 35896 14170 35902 14172
rect 35656 14118 35658 14170
rect 35838 14118 35840 14170
rect 35594 14116 35600 14118
rect 35656 14116 35680 14118
rect 35736 14116 35760 14118
rect 35816 14116 35840 14118
rect 35896 14116 35902 14118
rect 35594 14107 35902 14116
rect 27896 14068 27948 14074
rect 27896 14010 27948 14016
rect 27712 13932 27764 13938
rect 27712 13874 27764 13880
rect 27724 13530 27752 13874
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 27712 13524 27764 13530
rect 27712 13466 27764 13472
rect 27528 13320 27580 13326
rect 27528 13262 27580 13268
rect 28080 13320 28132 13326
rect 28080 13262 28132 13268
rect 27344 12980 27396 12986
rect 27344 12922 27396 12928
rect 26792 12844 26844 12850
rect 26792 12786 26844 12792
rect 26804 12434 26832 12786
rect 27540 12646 27568 13262
rect 27712 12776 27764 12782
rect 27712 12718 27764 12724
rect 27528 12640 27580 12646
rect 27528 12582 27580 12588
rect 26804 12406 26924 12434
rect 26896 12238 26924 12406
rect 26884 12232 26936 12238
rect 26884 12174 26936 12180
rect 26976 12232 27028 12238
rect 26976 12174 27028 12180
rect 27252 12232 27304 12238
rect 27252 12174 27304 12180
rect 26884 11756 26936 11762
rect 26988 11744 27016 12174
rect 26936 11716 27016 11744
rect 26884 11698 26936 11704
rect 26884 11348 26936 11354
rect 26884 11290 26936 11296
rect 26712 11070 26832 11098
rect 26424 11008 26476 11014
rect 26424 10950 26476 10956
rect 26700 11008 26752 11014
rect 26700 10950 26752 10956
rect 26436 10810 26464 10950
rect 26332 10804 26384 10810
rect 26332 10746 26384 10752
rect 26424 10804 26476 10810
rect 26424 10746 26476 10752
rect 26240 10736 26292 10742
rect 26240 10678 26292 10684
rect 26712 10470 26740 10950
rect 26700 10464 26752 10470
rect 26700 10406 26752 10412
rect 26240 10056 26292 10062
rect 26240 9998 26292 10004
rect 26252 9722 26280 9998
rect 26148 9716 26200 9722
rect 26148 9658 26200 9664
rect 26240 9716 26292 9722
rect 26240 9658 26292 9664
rect 26606 9616 26662 9625
rect 26148 9580 26200 9586
rect 26606 9551 26608 9560
rect 26148 9522 26200 9528
rect 26660 9551 26662 9560
rect 26608 9522 26660 9528
rect 26160 8838 26188 9522
rect 26700 9512 26752 9518
rect 26700 9454 26752 9460
rect 26516 9376 26568 9382
rect 26344 9336 26516 9364
rect 26148 8832 26200 8838
rect 26148 8774 26200 8780
rect 26344 8498 26372 9336
rect 26516 9318 26568 9324
rect 26712 9110 26740 9454
rect 26804 9178 26832 11070
rect 26896 11014 26924 11290
rect 26976 11144 27028 11150
rect 27264 11121 27292 12174
rect 27540 11694 27568 12582
rect 27724 12442 27752 12718
rect 27712 12436 27764 12442
rect 27712 12378 27764 12384
rect 28092 12306 28120 13262
rect 29920 13184 29972 13190
rect 29920 13126 29972 13132
rect 28816 12844 28868 12850
rect 28816 12786 28868 12792
rect 28080 12300 28132 12306
rect 28080 12242 28132 12248
rect 28172 12232 28224 12238
rect 28172 12174 28224 12180
rect 28724 12232 28776 12238
rect 28724 12174 28776 12180
rect 27620 12096 27672 12102
rect 27620 12038 27672 12044
rect 27528 11688 27580 11694
rect 27528 11630 27580 11636
rect 27344 11280 27396 11286
rect 27344 11222 27396 11228
rect 26976 11086 27028 11092
rect 27250 11112 27306 11121
rect 26884 11008 26936 11014
rect 26884 10950 26936 10956
rect 26988 10810 27016 11086
rect 27250 11047 27252 11056
rect 27304 11047 27306 11056
rect 27252 11018 27304 11024
rect 26976 10804 27028 10810
rect 26976 10746 27028 10752
rect 27264 10742 27292 11018
rect 27356 11014 27384 11222
rect 27344 11008 27396 11014
rect 27344 10950 27396 10956
rect 27356 10810 27384 10950
rect 27344 10804 27396 10810
rect 27344 10746 27396 10752
rect 27252 10736 27304 10742
rect 27252 10678 27304 10684
rect 27160 10464 27212 10470
rect 27160 10406 27212 10412
rect 26882 9616 26938 9625
rect 26938 9574 27016 9602
rect 26882 9551 26938 9560
rect 26884 9512 26936 9518
rect 26884 9454 26936 9460
rect 26792 9172 26844 9178
rect 26792 9114 26844 9120
rect 26700 9104 26752 9110
rect 26700 9046 26752 9052
rect 26332 8492 26384 8498
rect 26252 8452 26332 8480
rect 26056 7880 26108 7886
rect 26056 7822 26108 7828
rect 25872 7540 25924 7546
rect 25872 7482 25924 7488
rect 26252 6882 26280 8452
rect 26332 8434 26384 8440
rect 26424 8492 26476 8498
rect 26424 8434 26476 8440
rect 26332 7744 26384 7750
rect 26436 7732 26464 8434
rect 26896 8362 26924 9454
rect 26988 9382 27016 9574
rect 27068 9512 27120 9518
rect 27068 9454 27120 9460
rect 26976 9376 27028 9382
rect 26976 9318 27028 9324
rect 27080 8838 27108 9454
rect 27172 9382 27200 10406
rect 27540 10266 27568 11630
rect 27632 11558 27660 12038
rect 28184 11898 28212 12174
rect 28172 11892 28224 11898
rect 28172 11834 28224 11840
rect 27804 11688 27856 11694
rect 27804 11630 27856 11636
rect 27620 11552 27672 11558
rect 27620 11494 27672 11500
rect 27632 11150 27660 11494
rect 27816 11354 27844 11630
rect 27804 11348 27856 11354
rect 27804 11290 27856 11296
rect 27896 11348 27948 11354
rect 27896 11290 27948 11296
rect 27620 11144 27672 11150
rect 27620 11086 27672 11092
rect 27804 11144 27856 11150
rect 27804 11086 27856 11092
rect 27816 10810 27844 11086
rect 27908 10810 27936 11290
rect 27804 10804 27856 10810
rect 27804 10746 27856 10752
rect 27896 10804 27948 10810
rect 27896 10746 27948 10752
rect 27620 10600 27672 10606
rect 27620 10542 27672 10548
rect 27528 10260 27580 10266
rect 27528 10202 27580 10208
rect 27252 9988 27304 9994
rect 27252 9930 27304 9936
rect 27264 9654 27292 9930
rect 27632 9674 27660 10542
rect 28080 10056 28132 10062
rect 28080 9998 28132 10004
rect 27712 9920 27764 9926
rect 27712 9862 27764 9868
rect 27252 9648 27304 9654
rect 27252 9590 27304 9596
rect 27448 9646 27660 9674
rect 27724 9654 27752 9862
rect 27712 9648 27764 9654
rect 27448 9518 27476 9646
rect 27712 9590 27764 9596
rect 27436 9512 27488 9518
rect 27436 9454 27488 9460
rect 27344 9444 27396 9450
rect 27344 9386 27396 9392
rect 27160 9376 27212 9382
rect 27160 9318 27212 9324
rect 27356 9042 27384 9386
rect 27344 9036 27396 9042
rect 27344 8978 27396 8984
rect 27068 8832 27120 8838
rect 27068 8774 27120 8780
rect 27448 8634 27476 9454
rect 28092 9042 28120 9998
rect 28736 9994 28764 12174
rect 28828 11762 28856 12786
rect 29552 12776 29604 12782
rect 29552 12718 29604 12724
rect 29564 12374 29592 12718
rect 29552 12368 29604 12374
rect 29552 12310 29604 12316
rect 28816 11756 28868 11762
rect 28816 11698 28868 11704
rect 28828 10742 28856 11698
rect 29564 11354 29592 12310
rect 29736 12096 29788 12102
rect 29736 12038 29788 12044
rect 29644 11756 29696 11762
rect 29644 11698 29696 11704
rect 29552 11348 29604 11354
rect 29552 11290 29604 11296
rect 29564 11150 29592 11290
rect 29656 11150 29684 11698
rect 29748 11558 29776 12038
rect 29932 11626 29960 13126
rect 35594 13084 35902 13093
rect 35594 13082 35600 13084
rect 35656 13082 35680 13084
rect 35736 13082 35760 13084
rect 35816 13082 35840 13084
rect 35896 13082 35902 13084
rect 35656 13030 35658 13082
rect 35838 13030 35840 13082
rect 35594 13028 35600 13030
rect 35656 13028 35680 13030
rect 35736 13028 35760 13030
rect 35816 13028 35840 13030
rect 35896 13028 35902 13030
rect 35594 13019 35902 13028
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 35594 11996 35902 12005
rect 35594 11994 35600 11996
rect 35656 11994 35680 11996
rect 35736 11994 35760 11996
rect 35816 11994 35840 11996
rect 35896 11994 35902 11996
rect 35656 11942 35658 11994
rect 35838 11942 35840 11994
rect 35594 11940 35600 11942
rect 35656 11940 35680 11942
rect 35736 11940 35760 11942
rect 35816 11940 35840 11942
rect 35896 11940 35902 11942
rect 35594 11931 35902 11940
rect 29920 11620 29972 11626
rect 29920 11562 29972 11568
rect 38200 11620 38252 11626
rect 38200 11562 38252 11568
rect 29736 11552 29788 11558
rect 29736 11494 29788 11500
rect 29828 11552 29880 11558
rect 29828 11494 29880 11500
rect 29748 11150 29776 11494
rect 29840 11354 29868 11494
rect 29828 11348 29880 11354
rect 29828 11290 29880 11296
rect 29932 11218 29960 11562
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 29920 11212 29972 11218
rect 29920 11154 29972 11160
rect 29552 11144 29604 11150
rect 29552 11086 29604 11092
rect 29644 11144 29696 11150
rect 29644 11086 29696 11092
rect 29736 11144 29788 11150
rect 29736 11086 29788 11092
rect 29656 10810 29684 11086
rect 30012 11008 30064 11014
rect 30012 10950 30064 10956
rect 29644 10804 29696 10810
rect 29644 10746 29696 10752
rect 28816 10736 28868 10742
rect 28816 10678 28868 10684
rect 30024 10062 30052 10950
rect 35594 10908 35902 10917
rect 35594 10906 35600 10908
rect 35656 10906 35680 10908
rect 35736 10906 35760 10908
rect 35816 10906 35840 10908
rect 35896 10906 35902 10908
rect 35656 10854 35658 10906
rect 35838 10854 35840 10906
rect 35594 10852 35600 10854
rect 35656 10852 35680 10854
rect 35736 10852 35760 10854
rect 35816 10852 35840 10854
rect 35896 10852 35902 10854
rect 35594 10843 35902 10852
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 30012 10056 30064 10062
rect 30012 9998 30064 10004
rect 30104 10056 30156 10062
rect 30104 9998 30156 10004
rect 28172 9988 28224 9994
rect 28172 9930 28224 9936
rect 28632 9988 28684 9994
rect 28632 9930 28684 9936
rect 28724 9988 28776 9994
rect 28724 9930 28776 9936
rect 28184 9625 28212 9930
rect 28264 9648 28316 9654
rect 28170 9616 28226 9625
rect 28264 9590 28316 9596
rect 28170 9551 28226 9560
rect 28276 9178 28304 9590
rect 28448 9376 28500 9382
rect 28500 9336 28580 9364
rect 28448 9318 28500 9324
rect 28552 9178 28580 9336
rect 28644 9178 28672 9930
rect 30024 9178 30052 9998
rect 30116 9722 30144 9998
rect 35594 9820 35902 9829
rect 35594 9818 35600 9820
rect 35656 9818 35680 9820
rect 35736 9818 35760 9820
rect 35816 9818 35840 9820
rect 35896 9818 35902 9820
rect 35656 9766 35658 9818
rect 35838 9766 35840 9818
rect 35594 9764 35600 9766
rect 35656 9764 35680 9766
rect 35736 9764 35760 9766
rect 35816 9764 35840 9766
rect 35896 9764 35902 9766
rect 35594 9755 35902 9764
rect 30104 9716 30156 9722
rect 30104 9658 30156 9664
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 28264 9172 28316 9178
rect 28264 9114 28316 9120
rect 28540 9172 28592 9178
rect 28540 9114 28592 9120
rect 28632 9172 28684 9178
rect 28632 9114 28684 9120
rect 30012 9172 30064 9178
rect 30012 9114 30064 9120
rect 28080 9036 28132 9042
rect 28080 8978 28132 8984
rect 28172 8968 28224 8974
rect 28092 8916 28172 8922
rect 28092 8910 28224 8916
rect 28092 8894 28212 8910
rect 28092 8838 28120 8894
rect 27804 8832 27856 8838
rect 27804 8774 27856 8780
rect 27896 8832 27948 8838
rect 27896 8774 27948 8780
rect 28080 8832 28132 8838
rect 28080 8774 28132 8780
rect 27436 8628 27488 8634
rect 27436 8570 27488 8576
rect 26884 8356 26936 8362
rect 26884 8298 26936 8304
rect 27448 8090 27476 8570
rect 27816 8498 27844 8774
rect 27908 8566 27936 8774
rect 27896 8560 27948 8566
rect 27896 8502 27948 8508
rect 28092 8498 28120 8774
rect 28276 8566 28304 9114
rect 28552 8888 28580 9114
rect 29736 9104 29788 9110
rect 29736 9046 29788 9052
rect 28724 8900 28776 8906
rect 28552 8860 28724 8888
rect 28724 8842 28776 8848
rect 28264 8560 28316 8566
rect 28264 8502 28316 8508
rect 27528 8492 27580 8498
rect 27528 8434 27580 8440
rect 27620 8492 27672 8498
rect 27620 8434 27672 8440
rect 27804 8492 27856 8498
rect 27804 8434 27856 8440
rect 28080 8492 28132 8498
rect 28080 8434 28132 8440
rect 27068 8084 27120 8090
rect 27068 8026 27120 8032
rect 27436 8084 27488 8090
rect 27436 8026 27488 8032
rect 26384 7704 26464 7732
rect 26332 7686 26384 7692
rect 26344 6934 26372 7686
rect 26516 7404 26568 7410
rect 26516 7346 26568 7352
rect 26608 7404 26660 7410
rect 26608 7346 26660 7352
rect 26976 7404 27028 7410
rect 26976 7346 27028 7352
rect 26068 6854 26280 6882
rect 26332 6928 26384 6934
rect 26332 6870 26384 6876
rect 26068 6798 26096 6854
rect 26056 6792 26108 6798
rect 26056 6734 26108 6740
rect 26332 6792 26384 6798
rect 26332 6734 26384 6740
rect 26068 6662 26096 6734
rect 26056 6656 26108 6662
rect 26056 6598 26108 6604
rect 26344 6458 26372 6734
rect 26528 6730 26556 7346
rect 26620 6798 26648 7346
rect 26700 7200 26752 7206
rect 26700 7142 26752 7148
rect 26712 7002 26740 7142
rect 26700 6996 26752 7002
rect 26700 6938 26752 6944
rect 26608 6792 26660 6798
rect 26608 6734 26660 6740
rect 26516 6724 26568 6730
rect 26516 6666 26568 6672
rect 25780 6452 25832 6458
rect 25780 6394 25832 6400
rect 26332 6452 26384 6458
rect 26332 6394 26384 6400
rect 25792 6186 25820 6394
rect 25780 6180 25832 6186
rect 25780 6122 25832 6128
rect 25688 5908 25740 5914
rect 25688 5850 25740 5856
rect 25792 5710 25820 6122
rect 26528 6118 26556 6666
rect 26620 6322 26648 6734
rect 26608 6316 26660 6322
rect 26608 6258 26660 6264
rect 26240 6112 26292 6118
rect 26240 6054 26292 6060
rect 26516 6112 26568 6118
rect 26516 6054 26568 6060
rect 25780 5704 25832 5710
rect 25780 5646 25832 5652
rect 26252 5370 26280 6054
rect 26620 5914 26648 6258
rect 26608 5908 26660 5914
rect 26608 5850 26660 5856
rect 26516 5636 26568 5642
rect 26516 5578 26568 5584
rect 26528 5370 26556 5578
rect 26712 5574 26740 6938
rect 26988 6798 27016 7346
rect 26976 6792 27028 6798
rect 26976 6734 27028 6740
rect 26988 6662 27016 6734
rect 26976 6656 27028 6662
rect 26976 6598 27028 6604
rect 27080 5778 27108 8026
rect 27160 7336 27212 7342
rect 27160 7278 27212 7284
rect 27344 7336 27396 7342
rect 27344 7278 27396 7284
rect 27172 6934 27200 7278
rect 27356 7206 27384 7278
rect 27540 7274 27568 8434
rect 27632 7410 27660 8434
rect 28276 8090 28304 8502
rect 28632 8424 28684 8430
rect 28632 8366 28684 8372
rect 28356 8288 28408 8294
rect 28356 8230 28408 8236
rect 28448 8288 28500 8294
rect 28448 8230 28500 8236
rect 27988 8084 28040 8090
rect 27988 8026 28040 8032
rect 28264 8084 28316 8090
rect 28264 8026 28316 8032
rect 27804 7948 27856 7954
rect 27804 7890 27856 7896
rect 27620 7404 27672 7410
rect 27620 7346 27672 7352
rect 27816 7342 27844 7890
rect 27896 7812 27948 7818
rect 27896 7754 27948 7760
rect 27908 7478 27936 7754
rect 27896 7472 27948 7478
rect 27896 7414 27948 7420
rect 27908 7342 27936 7414
rect 27804 7336 27856 7342
rect 27804 7278 27856 7284
rect 27896 7336 27948 7342
rect 27896 7278 27948 7284
rect 27528 7268 27580 7274
rect 27528 7210 27580 7216
rect 27344 7200 27396 7206
rect 27344 7142 27396 7148
rect 27710 7168 27766 7177
rect 27710 7103 27766 7112
rect 27160 6928 27212 6934
rect 27160 6870 27212 6876
rect 27724 6798 27752 7103
rect 27816 7002 27844 7278
rect 28000 7018 28028 8026
rect 28368 7886 28396 8230
rect 28356 7880 28408 7886
rect 28356 7822 28408 7828
rect 28264 7404 28316 7410
rect 28264 7346 28316 7352
rect 28276 7177 28304 7346
rect 28368 7274 28396 7822
rect 28460 7750 28488 8230
rect 28644 7954 28672 8366
rect 28632 7948 28684 7954
rect 28632 7890 28684 7896
rect 28448 7744 28500 7750
rect 28448 7686 28500 7692
rect 28460 7410 28488 7686
rect 28448 7404 28500 7410
rect 28448 7346 28500 7352
rect 28356 7268 28408 7274
rect 28356 7210 28408 7216
rect 28262 7168 28318 7177
rect 28736 7154 28764 8842
rect 29552 8832 29604 8838
rect 29552 8774 29604 8780
rect 28908 8628 28960 8634
rect 28908 8570 28960 8576
rect 28920 7478 28948 8570
rect 29276 8084 29328 8090
rect 29276 8026 29328 8032
rect 29288 7478 29316 8026
rect 29564 7954 29592 8774
rect 29644 8560 29696 8566
rect 29644 8502 29696 8508
rect 29656 8090 29684 8502
rect 29644 8084 29696 8090
rect 29644 8026 29696 8032
rect 29748 7954 29776 9046
rect 35594 8732 35902 8741
rect 35594 8730 35600 8732
rect 35656 8730 35680 8732
rect 35736 8730 35760 8732
rect 35816 8730 35840 8732
rect 35896 8730 35902 8732
rect 35656 8678 35658 8730
rect 35838 8678 35840 8730
rect 35594 8676 35600 8678
rect 35656 8676 35680 8678
rect 35736 8676 35760 8678
rect 35816 8676 35840 8678
rect 35896 8676 35902 8678
rect 35594 8667 35902 8676
rect 38212 8634 38240 11562
rect 38200 8628 38252 8634
rect 38200 8570 38252 8576
rect 30012 8492 30064 8498
rect 30012 8434 30064 8440
rect 30196 8492 30248 8498
rect 30196 8434 30248 8440
rect 30564 8492 30616 8498
rect 30564 8434 30616 8440
rect 29828 8288 29880 8294
rect 29828 8230 29880 8236
rect 29552 7948 29604 7954
rect 29552 7890 29604 7896
rect 29736 7948 29788 7954
rect 29736 7890 29788 7896
rect 28908 7472 28960 7478
rect 28908 7414 28960 7420
rect 29092 7472 29144 7478
rect 29092 7414 29144 7420
rect 29276 7472 29328 7478
rect 29276 7414 29328 7420
rect 28318 7126 28764 7154
rect 28908 7200 28960 7206
rect 28908 7142 28960 7148
rect 28262 7103 28318 7112
rect 27804 6996 27856 7002
rect 27804 6938 27856 6944
rect 27908 6990 28028 7018
rect 28632 6996 28684 7002
rect 27436 6792 27488 6798
rect 27434 6760 27436 6769
rect 27620 6792 27672 6798
rect 27488 6760 27490 6769
rect 27620 6734 27672 6740
rect 27712 6792 27764 6798
rect 27712 6734 27764 6740
rect 27434 6695 27490 6704
rect 27436 6656 27488 6662
rect 27436 6598 27488 6604
rect 27448 6322 27476 6598
rect 27632 6458 27660 6734
rect 27620 6452 27672 6458
rect 27620 6394 27672 6400
rect 27436 6316 27488 6322
rect 27436 6258 27488 6264
rect 27160 6180 27212 6186
rect 27160 6122 27212 6128
rect 27068 5772 27120 5778
rect 27068 5714 27120 5720
rect 26700 5568 26752 5574
rect 26700 5510 26752 5516
rect 24400 5364 24452 5370
rect 24400 5306 24452 5312
rect 26240 5364 26292 5370
rect 26240 5306 26292 5312
rect 26516 5364 26568 5370
rect 26516 5306 26568 5312
rect 26424 5160 26476 5166
rect 26424 5102 26476 5108
rect 26436 4826 26464 5102
rect 26424 4820 26476 4826
rect 26424 4762 26476 4768
rect 27172 4622 27200 6122
rect 27448 4622 27476 6258
rect 27724 6186 27752 6734
rect 27908 6390 27936 6990
rect 28632 6938 28684 6944
rect 28446 6896 28502 6905
rect 28368 6854 28446 6882
rect 27986 6760 28042 6769
rect 27986 6695 28042 6704
rect 27896 6384 27948 6390
rect 27896 6326 27948 6332
rect 27712 6180 27764 6186
rect 27712 6122 27764 6128
rect 27908 5710 27936 6326
rect 28000 5914 28028 6695
rect 28368 6662 28396 6854
rect 28446 6831 28502 6840
rect 28448 6792 28500 6798
rect 28500 6752 28580 6780
rect 28644 6769 28672 6938
rect 28448 6734 28500 6740
rect 28356 6656 28408 6662
rect 28356 6598 28408 6604
rect 28448 6656 28500 6662
rect 28448 6598 28500 6604
rect 27988 5908 28040 5914
rect 27988 5850 28040 5856
rect 27896 5704 27948 5710
rect 27896 5646 27948 5652
rect 28000 5234 28028 5850
rect 28172 5568 28224 5574
rect 28172 5510 28224 5516
rect 28184 5370 28212 5510
rect 28172 5364 28224 5370
rect 28172 5306 28224 5312
rect 27988 5228 28040 5234
rect 27988 5170 28040 5176
rect 28368 4826 28396 6598
rect 28460 5914 28488 6598
rect 28552 6254 28580 6752
rect 28630 6760 28686 6769
rect 28736 6746 28764 7126
rect 28816 6996 28868 7002
rect 28816 6938 28868 6944
rect 28828 6905 28856 6938
rect 28814 6896 28870 6905
rect 28920 6866 28948 7142
rect 28814 6831 28870 6840
rect 28908 6860 28960 6866
rect 28908 6802 28960 6808
rect 28736 6730 28948 6746
rect 28736 6724 28960 6730
rect 28736 6718 28908 6724
rect 28630 6695 28686 6704
rect 28908 6666 28960 6672
rect 28816 6656 28868 6662
rect 28816 6598 28868 6604
rect 28828 6458 28856 6598
rect 29104 6458 29132 7414
rect 29748 7002 29776 7890
rect 29840 7410 29868 8230
rect 30024 7886 30052 8434
rect 30012 7880 30064 7886
rect 30012 7822 30064 7828
rect 29828 7404 29880 7410
rect 29828 7346 29880 7352
rect 30024 7002 30052 7822
rect 30208 7546 30236 8434
rect 30576 8090 30604 8434
rect 38844 8356 38896 8362
rect 38844 8298 38896 8304
rect 38856 8265 38884 8298
rect 38842 8256 38898 8265
rect 34934 8188 35242 8197
rect 38842 8191 38898 8200
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 30564 8084 30616 8090
rect 30564 8026 30616 8032
rect 30288 7880 30340 7886
rect 30288 7822 30340 7828
rect 30300 7546 30328 7822
rect 35594 7644 35902 7653
rect 35594 7642 35600 7644
rect 35656 7642 35680 7644
rect 35736 7642 35760 7644
rect 35816 7642 35840 7644
rect 35896 7642 35902 7644
rect 35656 7590 35658 7642
rect 35838 7590 35840 7642
rect 35594 7588 35600 7590
rect 35656 7588 35680 7590
rect 35736 7588 35760 7590
rect 35816 7588 35840 7590
rect 35896 7588 35902 7590
rect 35594 7579 35902 7588
rect 30196 7540 30248 7546
rect 30196 7482 30248 7488
rect 30288 7540 30340 7546
rect 30288 7482 30340 7488
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 29736 6996 29788 7002
rect 29736 6938 29788 6944
rect 30012 6996 30064 7002
rect 30012 6938 30064 6944
rect 35594 6556 35902 6565
rect 35594 6554 35600 6556
rect 35656 6554 35680 6556
rect 35736 6554 35760 6556
rect 35816 6554 35840 6556
rect 35896 6554 35902 6556
rect 35656 6502 35658 6554
rect 35838 6502 35840 6554
rect 35594 6500 35600 6502
rect 35656 6500 35680 6502
rect 35736 6500 35760 6502
rect 35816 6500 35840 6502
rect 35896 6500 35902 6502
rect 35594 6491 35902 6500
rect 28816 6452 28868 6458
rect 28816 6394 28868 6400
rect 29092 6452 29144 6458
rect 29092 6394 29144 6400
rect 28540 6248 28592 6254
rect 28540 6190 28592 6196
rect 28448 5908 28500 5914
rect 28448 5850 28500 5856
rect 28828 5710 28856 6394
rect 29092 6248 29144 6254
rect 29092 6190 29144 6196
rect 29104 5914 29132 6190
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 29092 5908 29144 5914
rect 29092 5850 29144 5856
rect 28816 5704 28868 5710
rect 28816 5646 28868 5652
rect 29092 5568 29144 5574
rect 29092 5510 29144 5516
rect 29104 5370 29132 5510
rect 35594 5468 35902 5477
rect 35594 5466 35600 5468
rect 35656 5466 35680 5468
rect 35736 5466 35760 5468
rect 35816 5466 35840 5468
rect 35896 5466 35902 5468
rect 35656 5414 35658 5466
rect 35838 5414 35840 5466
rect 35594 5412 35600 5414
rect 35656 5412 35680 5414
rect 35736 5412 35760 5414
rect 35816 5412 35840 5414
rect 35896 5412 35902 5414
rect 35594 5403 35902 5412
rect 29092 5364 29144 5370
rect 29092 5306 29144 5312
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 28356 4820 28408 4826
rect 28356 4762 28408 4768
rect 27160 4616 27212 4622
rect 27160 4558 27212 4564
rect 27436 4616 27488 4622
rect 27436 4558 27488 4564
rect 35594 4380 35902 4389
rect 35594 4378 35600 4380
rect 35656 4378 35680 4380
rect 35736 4378 35760 4380
rect 35816 4378 35840 4380
rect 35896 4378 35902 4380
rect 35656 4326 35658 4378
rect 35838 4326 35840 4378
rect 35594 4324 35600 4326
rect 35656 4324 35680 4326
rect 35736 4324 35760 4326
rect 35816 4324 35840 4326
rect 35896 4324 35902 4326
rect 35594 4315 35902 4324
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35594 3292 35902 3301
rect 35594 3290 35600 3292
rect 35656 3290 35680 3292
rect 35736 3290 35760 3292
rect 35816 3290 35840 3292
rect 35896 3290 35902 3292
rect 35656 3238 35658 3290
rect 35838 3238 35840 3290
rect 35594 3236 35600 3238
rect 35656 3236 35680 3238
rect 35736 3236 35760 3238
rect 35816 3236 35840 3238
rect 35896 3236 35902 3238
rect 35594 3227 35902 3236
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 24216 2644 24268 2650
rect 24216 2586 24268 2592
rect 23848 2440 23900 2446
rect 23848 2382 23900 2388
rect 22100 2372 22152 2378
rect 22100 2314 22152 2320
rect 18696 2304 18748 2310
rect 18696 2246 18748 2252
rect 22008 2304 22060 2310
rect 22008 2246 22060 2252
rect 11624 1142 11836 1170
rect 11624 800 11652 1142
rect 23860 800 23888 2382
rect 35440 2304 35492 2310
rect 35440 2246 35492 2252
rect 35452 800 35480 2246
rect 35594 2204 35902 2213
rect 35594 2202 35600 2204
rect 35656 2202 35680 2204
rect 35736 2202 35760 2204
rect 35816 2202 35840 2204
rect 35896 2202 35902 2204
rect 35656 2150 35658 2202
rect 35838 2150 35840 2202
rect 35594 2148 35600 2150
rect 35656 2148 35680 2150
rect 35736 2148 35760 2150
rect 35816 2148 35840 2150
rect 35896 2148 35902 2150
rect 35594 2139 35902 2148
rect 18 0 74 800
rect 11610 0 11666 800
rect 23846 0 23902 800
rect 35438 0 35494 800
<< via2 >>
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 938 37460 994 37496
rect 938 37440 940 37460
rect 940 37440 992 37460
rect 992 37440 994 37460
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 938 25220 994 25256
rect 938 25200 940 25220
rect 940 25200 992 25220
rect 992 25200 994 25220
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 1398 12280 1454 12336
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 20442 11892 20498 11928
rect 20442 11872 20444 11892
rect 20444 11872 20496 11892
rect 20496 11872 20498 11892
rect 35600 37018 35656 37020
rect 35680 37018 35736 37020
rect 35760 37018 35816 37020
rect 35840 37018 35896 37020
rect 35600 36966 35646 37018
rect 35646 36966 35656 37018
rect 35680 36966 35710 37018
rect 35710 36966 35722 37018
rect 35722 36966 35736 37018
rect 35760 36966 35774 37018
rect 35774 36966 35786 37018
rect 35786 36966 35816 37018
rect 35840 36966 35850 37018
rect 35850 36966 35896 37018
rect 35600 36964 35656 36966
rect 35680 36964 35736 36966
rect 35760 36964 35816 36966
rect 35840 36964 35896 36966
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 35600 35930 35656 35932
rect 35680 35930 35736 35932
rect 35760 35930 35816 35932
rect 35840 35930 35896 35932
rect 35600 35878 35646 35930
rect 35646 35878 35656 35930
rect 35680 35878 35710 35930
rect 35710 35878 35722 35930
rect 35722 35878 35736 35930
rect 35760 35878 35774 35930
rect 35774 35878 35786 35930
rect 35786 35878 35816 35930
rect 35840 35878 35850 35930
rect 35850 35878 35896 35930
rect 35600 35876 35656 35878
rect 35680 35876 35736 35878
rect 35760 35876 35816 35878
rect 35840 35876 35896 35878
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 35600 34842 35656 34844
rect 35680 34842 35736 34844
rect 35760 34842 35816 34844
rect 35840 34842 35896 34844
rect 35600 34790 35646 34842
rect 35646 34790 35656 34842
rect 35680 34790 35710 34842
rect 35710 34790 35722 34842
rect 35722 34790 35736 34842
rect 35760 34790 35774 34842
rect 35774 34790 35786 34842
rect 35786 34790 35816 34842
rect 35840 34790 35850 34842
rect 35850 34790 35896 34842
rect 35600 34788 35656 34790
rect 35680 34788 35736 34790
rect 35760 34788 35816 34790
rect 35840 34788 35896 34790
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 35600 33754 35656 33756
rect 35680 33754 35736 33756
rect 35760 33754 35816 33756
rect 35840 33754 35896 33756
rect 35600 33702 35646 33754
rect 35646 33702 35656 33754
rect 35680 33702 35710 33754
rect 35710 33702 35722 33754
rect 35722 33702 35736 33754
rect 35760 33702 35774 33754
rect 35774 33702 35786 33754
rect 35786 33702 35816 33754
rect 35840 33702 35850 33754
rect 35850 33702 35896 33754
rect 35600 33700 35656 33702
rect 35680 33700 35736 33702
rect 35760 33700 35816 33702
rect 35840 33700 35896 33702
rect 38842 33360 38898 33416
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 35600 32666 35656 32668
rect 35680 32666 35736 32668
rect 35760 32666 35816 32668
rect 35840 32666 35896 32668
rect 35600 32614 35646 32666
rect 35646 32614 35656 32666
rect 35680 32614 35710 32666
rect 35710 32614 35722 32666
rect 35722 32614 35736 32666
rect 35760 32614 35774 32666
rect 35774 32614 35786 32666
rect 35786 32614 35816 32666
rect 35840 32614 35850 32666
rect 35850 32614 35896 32666
rect 35600 32612 35656 32614
rect 35680 32612 35736 32614
rect 35760 32612 35816 32614
rect 35840 32612 35896 32614
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 35600 31578 35656 31580
rect 35680 31578 35736 31580
rect 35760 31578 35816 31580
rect 35840 31578 35896 31580
rect 35600 31526 35646 31578
rect 35646 31526 35656 31578
rect 35680 31526 35710 31578
rect 35710 31526 35722 31578
rect 35722 31526 35736 31578
rect 35760 31526 35774 31578
rect 35774 31526 35786 31578
rect 35786 31526 35816 31578
rect 35840 31526 35850 31578
rect 35850 31526 35896 31578
rect 35600 31524 35656 31526
rect 35680 31524 35736 31526
rect 35760 31524 35816 31526
rect 35840 31524 35896 31526
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 35600 30490 35656 30492
rect 35680 30490 35736 30492
rect 35760 30490 35816 30492
rect 35840 30490 35896 30492
rect 35600 30438 35646 30490
rect 35646 30438 35656 30490
rect 35680 30438 35710 30490
rect 35710 30438 35722 30490
rect 35722 30438 35736 30490
rect 35760 30438 35774 30490
rect 35774 30438 35786 30490
rect 35786 30438 35816 30490
rect 35840 30438 35850 30490
rect 35850 30438 35896 30490
rect 35600 30436 35656 30438
rect 35680 30436 35736 30438
rect 35760 30436 35816 30438
rect 35840 30436 35896 30438
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 35600 29402 35656 29404
rect 35680 29402 35736 29404
rect 35760 29402 35816 29404
rect 35840 29402 35896 29404
rect 35600 29350 35646 29402
rect 35646 29350 35656 29402
rect 35680 29350 35710 29402
rect 35710 29350 35722 29402
rect 35722 29350 35736 29402
rect 35760 29350 35774 29402
rect 35774 29350 35786 29402
rect 35786 29350 35816 29402
rect 35840 29350 35850 29402
rect 35850 29350 35896 29402
rect 35600 29348 35656 29350
rect 35680 29348 35736 29350
rect 35760 29348 35816 29350
rect 35840 29348 35896 29350
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 35600 28314 35656 28316
rect 35680 28314 35736 28316
rect 35760 28314 35816 28316
rect 35840 28314 35896 28316
rect 35600 28262 35646 28314
rect 35646 28262 35656 28314
rect 35680 28262 35710 28314
rect 35710 28262 35722 28314
rect 35722 28262 35736 28314
rect 35760 28262 35774 28314
rect 35774 28262 35786 28314
rect 35786 28262 35816 28314
rect 35840 28262 35850 28314
rect 35850 28262 35896 28314
rect 35600 28260 35656 28262
rect 35680 28260 35736 28262
rect 35760 28260 35816 28262
rect 35840 28260 35896 28262
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 35600 27226 35656 27228
rect 35680 27226 35736 27228
rect 35760 27226 35816 27228
rect 35840 27226 35896 27228
rect 35600 27174 35646 27226
rect 35646 27174 35656 27226
rect 35680 27174 35710 27226
rect 35710 27174 35722 27226
rect 35722 27174 35736 27226
rect 35760 27174 35774 27226
rect 35774 27174 35786 27226
rect 35786 27174 35816 27226
rect 35840 27174 35850 27226
rect 35850 27174 35896 27226
rect 35600 27172 35656 27174
rect 35680 27172 35736 27174
rect 35760 27172 35816 27174
rect 35840 27172 35896 27174
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 35600 26138 35656 26140
rect 35680 26138 35736 26140
rect 35760 26138 35816 26140
rect 35840 26138 35896 26140
rect 35600 26086 35646 26138
rect 35646 26086 35656 26138
rect 35680 26086 35710 26138
rect 35710 26086 35722 26138
rect 35722 26086 35736 26138
rect 35760 26086 35774 26138
rect 35774 26086 35786 26138
rect 35786 26086 35816 26138
rect 35840 26086 35850 26138
rect 35850 26086 35896 26138
rect 35600 26084 35656 26086
rect 35680 26084 35736 26086
rect 35760 26084 35816 26086
rect 35840 26084 35896 26086
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 35600 25050 35656 25052
rect 35680 25050 35736 25052
rect 35760 25050 35816 25052
rect 35840 25050 35896 25052
rect 35600 24998 35646 25050
rect 35646 24998 35656 25050
rect 35680 24998 35710 25050
rect 35710 24998 35722 25050
rect 35722 24998 35736 25050
rect 35760 24998 35774 25050
rect 35774 24998 35786 25050
rect 35786 24998 35816 25050
rect 35840 24998 35850 25050
rect 35850 24998 35896 25050
rect 35600 24996 35656 24998
rect 35680 24996 35736 24998
rect 35760 24996 35816 24998
rect 35840 24996 35896 24998
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 35600 23962 35656 23964
rect 35680 23962 35736 23964
rect 35760 23962 35816 23964
rect 35840 23962 35896 23964
rect 35600 23910 35646 23962
rect 35646 23910 35656 23962
rect 35680 23910 35710 23962
rect 35710 23910 35722 23962
rect 35722 23910 35736 23962
rect 35760 23910 35774 23962
rect 35774 23910 35786 23962
rect 35786 23910 35816 23962
rect 35840 23910 35850 23962
rect 35850 23910 35896 23962
rect 35600 23908 35656 23910
rect 35680 23908 35736 23910
rect 35760 23908 35816 23910
rect 35840 23908 35896 23910
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 35600 22874 35656 22876
rect 35680 22874 35736 22876
rect 35760 22874 35816 22876
rect 35840 22874 35896 22876
rect 35600 22822 35646 22874
rect 35646 22822 35656 22874
rect 35680 22822 35710 22874
rect 35710 22822 35722 22874
rect 35722 22822 35736 22874
rect 35760 22822 35774 22874
rect 35774 22822 35786 22874
rect 35786 22822 35816 22874
rect 35840 22822 35850 22874
rect 35850 22822 35896 22874
rect 35600 22820 35656 22822
rect 35680 22820 35736 22822
rect 35760 22820 35816 22822
rect 35840 22820 35896 22822
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 35600 21786 35656 21788
rect 35680 21786 35736 21788
rect 35760 21786 35816 21788
rect 35840 21786 35896 21788
rect 35600 21734 35646 21786
rect 35646 21734 35656 21786
rect 35680 21734 35710 21786
rect 35710 21734 35722 21786
rect 35722 21734 35736 21786
rect 35760 21734 35774 21786
rect 35774 21734 35786 21786
rect 35786 21734 35816 21786
rect 35840 21734 35850 21786
rect 35850 21734 35896 21786
rect 35600 21732 35656 21734
rect 35680 21732 35736 21734
rect 35760 21732 35816 21734
rect 35840 21732 35896 21734
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 35600 20698 35656 20700
rect 35680 20698 35736 20700
rect 35760 20698 35816 20700
rect 35840 20698 35896 20700
rect 35600 20646 35646 20698
rect 35646 20646 35656 20698
rect 35680 20646 35710 20698
rect 35710 20646 35722 20698
rect 35722 20646 35736 20698
rect 35760 20646 35774 20698
rect 35774 20646 35786 20698
rect 35786 20646 35816 20698
rect 35840 20646 35850 20698
rect 35850 20646 35896 20698
rect 35600 20644 35656 20646
rect 35680 20644 35736 20646
rect 35760 20644 35816 20646
rect 35840 20644 35896 20646
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 35600 19610 35656 19612
rect 35680 19610 35736 19612
rect 35760 19610 35816 19612
rect 35840 19610 35896 19612
rect 35600 19558 35646 19610
rect 35646 19558 35656 19610
rect 35680 19558 35710 19610
rect 35710 19558 35722 19610
rect 35722 19558 35736 19610
rect 35760 19558 35774 19610
rect 35774 19558 35786 19610
rect 35786 19558 35816 19610
rect 35840 19558 35850 19610
rect 35850 19558 35896 19610
rect 35600 19556 35656 19558
rect 35680 19556 35736 19558
rect 35760 19556 35816 19558
rect 35840 19556 35896 19558
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 35600 18522 35656 18524
rect 35680 18522 35736 18524
rect 35760 18522 35816 18524
rect 35840 18522 35896 18524
rect 35600 18470 35646 18522
rect 35646 18470 35656 18522
rect 35680 18470 35710 18522
rect 35710 18470 35722 18522
rect 35722 18470 35736 18522
rect 35760 18470 35774 18522
rect 35774 18470 35786 18522
rect 35786 18470 35816 18522
rect 35840 18470 35850 18522
rect 35850 18470 35896 18522
rect 35600 18468 35656 18470
rect 35680 18468 35736 18470
rect 35760 18468 35816 18470
rect 35840 18468 35896 18470
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 35600 17434 35656 17436
rect 35680 17434 35736 17436
rect 35760 17434 35816 17436
rect 35840 17434 35896 17436
rect 35600 17382 35646 17434
rect 35646 17382 35656 17434
rect 35680 17382 35710 17434
rect 35710 17382 35722 17434
rect 35722 17382 35736 17434
rect 35760 17382 35774 17434
rect 35774 17382 35786 17434
rect 35786 17382 35816 17434
rect 35840 17382 35850 17434
rect 35850 17382 35896 17434
rect 35600 17380 35656 17382
rect 35680 17380 35736 17382
rect 35760 17380 35816 17382
rect 35840 17380 35896 17382
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 35600 16346 35656 16348
rect 35680 16346 35736 16348
rect 35760 16346 35816 16348
rect 35840 16346 35896 16348
rect 35600 16294 35646 16346
rect 35646 16294 35656 16346
rect 35680 16294 35710 16346
rect 35710 16294 35722 16346
rect 35722 16294 35736 16346
rect 35760 16294 35774 16346
rect 35774 16294 35786 16346
rect 35786 16294 35816 16346
rect 35840 16294 35850 16346
rect 35850 16294 35896 16346
rect 35600 16292 35656 16294
rect 35680 16292 35736 16294
rect 35760 16292 35816 16294
rect 35840 16292 35896 16294
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 35600 15258 35656 15260
rect 35680 15258 35736 15260
rect 35760 15258 35816 15260
rect 35840 15258 35896 15260
rect 35600 15206 35646 15258
rect 35646 15206 35656 15258
rect 35680 15206 35710 15258
rect 35710 15206 35722 15258
rect 35722 15206 35736 15258
rect 35760 15206 35774 15258
rect 35774 15206 35786 15258
rect 35786 15206 35816 15258
rect 35840 15206 35850 15258
rect 35850 15206 35896 15258
rect 35600 15204 35656 15206
rect 35680 15204 35736 15206
rect 35760 15204 35816 15206
rect 35840 15204 35896 15206
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 24674 11872 24730 11928
rect 25410 11092 25412 11112
rect 25412 11092 25464 11112
rect 25464 11092 25466 11112
rect 25410 11056 25466 11092
rect 25962 9560 26018 9616
rect 26238 11056 26294 11112
rect 26238 10920 26294 10976
rect 35600 14170 35656 14172
rect 35680 14170 35736 14172
rect 35760 14170 35816 14172
rect 35840 14170 35896 14172
rect 35600 14118 35646 14170
rect 35646 14118 35656 14170
rect 35680 14118 35710 14170
rect 35710 14118 35722 14170
rect 35722 14118 35736 14170
rect 35760 14118 35774 14170
rect 35774 14118 35786 14170
rect 35786 14118 35816 14170
rect 35840 14118 35850 14170
rect 35850 14118 35896 14170
rect 35600 14116 35656 14118
rect 35680 14116 35736 14118
rect 35760 14116 35816 14118
rect 35840 14116 35896 14118
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 26606 9580 26662 9616
rect 26606 9560 26608 9580
rect 26608 9560 26660 9580
rect 26660 9560 26662 9580
rect 27250 11076 27306 11112
rect 27250 11056 27252 11076
rect 27252 11056 27304 11076
rect 27304 11056 27306 11076
rect 26882 9560 26938 9616
rect 35600 13082 35656 13084
rect 35680 13082 35736 13084
rect 35760 13082 35816 13084
rect 35840 13082 35896 13084
rect 35600 13030 35646 13082
rect 35646 13030 35656 13082
rect 35680 13030 35710 13082
rect 35710 13030 35722 13082
rect 35722 13030 35736 13082
rect 35760 13030 35774 13082
rect 35774 13030 35786 13082
rect 35786 13030 35816 13082
rect 35840 13030 35850 13082
rect 35850 13030 35896 13082
rect 35600 13028 35656 13030
rect 35680 13028 35736 13030
rect 35760 13028 35816 13030
rect 35840 13028 35896 13030
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 35600 11994 35656 11996
rect 35680 11994 35736 11996
rect 35760 11994 35816 11996
rect 35840 11994 35896 11996
rect 35600 11942 35646 11994
rect 35646 11942 35656 11994
rect 35680 11942 35710 11994
rect 35710 11942 35722 11994
rect 35722 11942 35736 11994
rect 35760 11942 35774 11994
rect 35774 11942 35786 11994
rect 35786 11942 35816 11994
rect 35840 11942 35850 11994
rect 35850 11942 35896 11994
rect 35600 11940 35656 11942
rect 35680 11940 35736 11942
rect 35760 11940 35816 11942
rect 35840 11940 35896 11942
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 35600 10906 35656 10908
rect 35680 10906 35736 10908
rect 35760 10906 35816 10908
rect 35840 10906 35896 10908
rect 35600 10854 35646 10906
rect 35646 10854 35656 10906
rect 35680 10854 35710 10906
rect 35710 10854 35722 10906
rect 35722 10854 35736 10906
rect 35760 10854 35774 10906
rect 35774 10854 35786 10906
rect 35786 10854 35816 10906
rect 35840 10854 35850 10906
rect 35850 10854 35896 10906
rect 35600 10852 35656 10854
rect 35680 10852 35736 10854
rect 35760 10852 35816 10854
rect 35840 10852 35896 10854
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 28170 9560 28226 9616
rect 35600 9818 35656 9820
rect 35680 9818 35736 9820
rect 35760 9818 35816 9820
rect 35840 9818 35896 9820
rect 35600 9766 35646 9818
rect 35646 9766 35656 9818
rect 35680 9766 35710 9818
rect 35710 9766 35722 9818
rect 35722 9766 35736 9818
rect 35760 9766 35774 9818
rect 35774 9766 35786 9818
rect 35786 9766 35816 9818
rect 35840 9766 35850 9818
rect 35850 9766 35896 9818
rect 35600 9764 35656 9766
rect 35680 9764 35736 9766
rect 35760 9764 35816 9766
rect 35840 9764 35896 9766
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 27710 7112 27766 7168
rect 28262 7112 28318 7168
rect 35600 8730 35656 8732
rect 35680 8730 35736 8732
rect 35760 8730 35816 8732
rect 35840 8730 35896 8732
rect 35600 8678 35646 8730
rect 35646 8678 35656 8730
rect 35680 8678 35710 8730
rect 35710 8678 35722 8730
rect 35722 8678 35736 8730
rect 35760 8678 35774 8730
rect 35774 8678 35786 8730
rect 35786 8678 35816 8730
rect 35840 8678 35850 8730
rect 35850 8678 35896 8730
rect 35600 8676 35656 8678
rect 35680 8676 35736 8678
rect 35760 8676 35816 8678
rect 35840 8676 35896 8678
rect 27434 6740 27436 6760
rect 27436 6740 27488 6760
rect 27488 6740 27490 6760
rect 27434 6704 27490 6740
rect 27986 6704 28042 6760
rect 28446 6840 28502 6896
rect 28630 6704 28686 6760
rect 28814 6840 28870 6896
rect 38842 8200 38898 8256
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 35600 7642 35656 7644
rect 35680 7642 35736 7644
rect 35760 7642 35816 7644
rect 35840 7642 35896 7644
rect 35600 7590 35646 7642
rect 35646 7590 35656 7642
rect 35680 7590 35710 7642
rect 35710 7590 35722 7642
rect 35722 7590 35736 7642
rect 35760 7590 35774 7642
rect 35774 7590 35786 7642
rect 35786 7590 35816 7642
rect 35840 7590 35850 7642
rect 35850 7590 35896 7642
rect 35600 7588 35656 7590
rect 35680 7588 35736 7590
rect 35760 7588 35816 7590
rect 35840 7588 35896 7590
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 35600 6554 35656 6556
rect 35680 6554 35736 6556
rect 35760 6554 35816 6556
rect 35840 6554 35896 6556
rect 35600 6502 35646 6554
rect 35646 6502 35656 6554
rect 35680 6502 35710 6554
rect 35710 6502 35722 6554
rect 35722 6502 35736 6554
rect 35760 6502 35774 6554
rect 35774 6502 35786 6554
rect 35786 6502 35816 6554
rect 35840 6502 35850 6554
rect 35850 6502 35896 6554
rect 35600 6500 35656 6502
rect 35680 6500 35736 6502
rect 35760 6500 35816 6502
rect 35840 6500 35896 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 35600 5466 35656 5468
rect 35680 5466 35736 5468
rect 35760 5466 35816 5468
rect 35840 5466 35896 5468
rect 35600 5414 35646 5466
rect 35646 5414 35656 5466
rect 35680 5414 35710 5466
rect 35710 5414 35722 5466
rect 35722 5414 35736 5466
rect 35760 5414 35774 5466
rect 35774 5414 35786 5466
rect 35786 5414 35816 5466
rect 35840 5414 35850 5466
rect 35850 5414 35896 5466
rect 35600 5412 35656 5414
rect 35680 5412 35736 5414
rect 35760 5412 35816 5414
rect 35840 5412 35896 5414
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 35600 4378 35656 4380
rect 35680 4378 35736 4380
rect 35760 4378 35816 4380
rect 35840 4378 35896 4380
rect 35600 4326 35646 4378
rect 35646 4326 35656 4378
rect 35680 4326 35710 4378
rect 35710 4326 35722 4378
rect 35722 4326 35736 4378
rect 35760 4326 35774 4378
rect 35774 4326 35786 4378
rect 35786 4326 35816 4378
rect 35840 4326 35850 4378
rect 35850 4326 35896 4378
rect 35600 4324 35656 4326
rect 35680 4324 35736 4326
rect 35760 4324 35816 4326
rect 35840 4324 35896 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 35600 3290 35656 3292
rect 35680 3290 35736 3292
rect 35760 3290 35816 3292
rect 35840 3290 35896 3292
rect 35600 3238 35646 3290
rect 35646 3238 35656 3290
rect 35680 3238 35710 3290
rect 35710 3238 35722 3290
rect 35722 3238 35736 3290
rect 35760 3238 35774 3290
rect 35774 3238 35786 3290
rect 35786 3238 35816 3290
rect 35840 3238 35850 3290
rect 35850 3238 35896 3290
rect 35600 3236 35656 3238
rect 35680 3236 35736 3238
rect 35760 3236 35816 3238
rect 35840 3236 35896 3238
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35600 2202 35656 2204
rect 35680 2202 35736 2204
rect 35760 2202 35816 2204
rect 35840 2202 35896 2204
rect 35600 2150 35646 2202
rect 35646 2150 35656 2202
rect 35680 2150 35710 2202
rect 35710 2150 35722 2202
rect 35722 2150 35736 2202
rect 35760 2150 35774 2202
rect 35774 2150 35786 2202
rect 35786 2150 35816 2202
rect 35840 2150 35850 2202
rect 35850 2150 35896 2202
rect 35600 2148 35656 2150
rect 35680 2148 35736 2150
rect 35760 2148 35816 2150
rect 35840 2148 35896 2150
<< metal3 >>
rect 4210 37568 4526 37569
rect 0 37498 800 37528
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 933 37498 999 37501
rect 0 37496 999 37498
rect 0 37440 938 37496
rect 994 37440 999 37496
rect 0 37438 999 37440
rect 0 37408 800 37438
rect 933 37435 999 37438
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 35590 37024 35906 37025
rect 35590 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35906 37024
rect 35590 36959 35906 36960
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 35590 35936 35906 35937
rect 35590 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35906 35936
rect 35590 35871 35906 35872
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 4870 34848 5186 34849
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 35590 34848 35906 34849
rect 35590 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35906 34848
rect 35590 34783 35906 34784
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 35590 33760 35906 33761
rect 35590 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35906 33760
rect 35590 33695 35906 33696
rect 38837 33418 38903 33421
rect 39200 33418 40000 33448
rect 38837 33416 40000 33418
rect 38837 33360 38842 33416
rect 38898 33360 40000 33416
rect 38837 33358 40000 33360
rect 38837 33355 38903 33358
rect 39200 33328 40000 33358
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 35590 32672 35906 32673
rect 35590 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35906 32672
rect 35590 32607 35906 32608
rect 4210 32128 4526 32129
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 35590 31584 35906 31585
rect 35590 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35906 31584
rect 35590 31519 35906 31520
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 35590 30496 35906 30497
rect 35590 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35906 30496
rect 35590 30431 35906 30432
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 35590 29408 35906 29409
rect 35590 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35906 29408
rect 35590 29343 35906 29344
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 35590 28320 35906 28321
rect 35590 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35906 28320
rect 35590 28255 35906 28256
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 35590 27232 35906 27233
rect 35590 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35906 27232
rect 35590 27167 35906 27168
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 35590 26144 35906 26145
rect 35590 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35906 26144
rect 35590 26079 35906 26080
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 0 25258 800 25288
rect 933 25258 999 25261
rect 0 25256 999 25258
rect 0 25200 938 25256
rect 994 25200 999 25256
rect 0 25198 999 25200
rect 0 25168 800 25198
rect 933 25195 999 25198
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 35590 25056 35906 25057
rect 35590 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35906 25056
rect 35590 24991 35906 24992
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 35590 23968 35906 23969
rect 35590 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35906 23968
rect 35590 23903 35906 23904
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 35590 22880 35906 22881
rect 35590 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35906 22880
rect 35590 22815 35906 22816
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 35590 21792 35906 21793
rect 35590 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35906 21792
rect 35590 21727 35906 21728
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 39200 21178 40000 21208
rect 35850 21118 40000 21178
rect 34646 20980 34652 21044
rect 34716 21042 34722 21044
rect 35850 21042 35910 21118
rect 39200 21088 40000 21118
rect 34716 20982 35910 21042
rect 34716 20980 34722 20982
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 35590 20704 35906 20705
rect 35590 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35906 20704
rect 35590 20639 35906 20640
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 35590 19616 35906 19617
rect 35590 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35906 19616
rect 35590 19551 35906 19552
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 4870 18528 5186 18529
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 35590 18528 35906 18529
rect 35590 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35906 18528
rect 35590 18463 35906 18464
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 35590 17440 35906 17441
rect 35590 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35906 17440
rect 35590 17375 35906 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 35590 16352 35906 16353
rect 35590 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35906 16352
rect 35590 16287 35906 16288
rect 4210 15808 4526 15809
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 35590 15264 35906 15265
rect 35590 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35906 15264
rect 35590 15199 35906 15200
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 35590 14176 35906 14177
rect 35590 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35906 14176
rect 35590 14111 35906 14112
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 34930 13567 35246 13568
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 35590 13088 35906 13089
rect 35590 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35906 13088
rect 35590 13023 35906 13024
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 0 12338 800 12368
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 0 12248 800 12278
rect 1393 12275 1459 12278
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 35590 12000 35906 12001
rect 35590 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35906 12000
rect 35590 11935 35906 11936
rect 20437 11930 20503 11933
rect 24669 11930 24735 11933
rect 20437 11928 24735 11930
rect 20437 11872 20442 11928
rect 20498 11872 24674 11928
rect 24730 11872 24735 11928
rect 20437 11870 24735 11872
rect 20437 11867 20503 11870
rect 24669 11867 24735 11870
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 25405 11114 25471 11117
rect 26233 11114 26299 11117
rect 27245 11114 27311 11117
rect 25405 11112 27311 11114
rect 25405 11056 25410 11112
rect 25466 11056 26238 11112
rect 26294 11056 27250 11112
rect 27306 11056 27311 11112
rect 25405 11054 27311 11056
rect 25405 11051 25471 11054
rect 26233 11051 26299 11054
rect 27245 11051 27311 11054
rect 26233 10978 26299 10981
rect 34646 10978 34652 10980
rect 26233 10976 34652 10978
rect 26233 10920 26238 10976
rect 26294 10920 34652 10976
rect 26233 10918 34652 10920
rect 26233 10915 26299 10918
rect 34646 10916 34652 10918
rect 34716 10916 34722 10980
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 35590 10912 35906 10913
rect 35590 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35906 10912
rect 35590 10847 35906 10848
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 35590 9824 35906 9825
rect 35590 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35906 9824
rect 35590 9759 35906 9760
rect 25957 9618 26023 9621
rect 26601 9618 26667 9621
rect 25957 9616 26667 9618
rect 25957 9560 25962 9616
rect 26018 9560 26606 9616
rect 26662 9560 26667 9616
rect 25957 9558 26667 9560
rect 25957 9555 26023 9558
rect 26601 9555 26667 9558
rect 26877 9618 26943 9621
rect 28165 9618 28231 9621
rect 26877 9616 28231 9618
rect 26877 9560 26882 9616
rect 26938 9560 28170 9616
rect 28226 9560 28231 9616
rect 26877 9558 28231 9560
rect 26877 9555 26943 9558
rect 28165 9555 28231 9558
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 35590 8736 35906 8737
rect 35590 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35906 8736
rect 35590 8671 35906 8672
rect 38837 8258 38903 8261
rect 39200 8258 40000 8288
rect 38837 8256 40000 8258
rect 38837 8200 38842 8256
rect 38898 8200 40000 8256
rect 38837 8198 40000 8200
rect 38837 8195 38903 8198
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 39200 8168 40000 8198
rect 34930 8127 35246 8128
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 35590 7648 35906 7649
rect 35590 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35906 7648
rect 35590 7583 35906 7584
rect 27705 7170 27771 7173
rect 28257 7170 28323 7173
rect 27705 7168 28323 7170
rect 27705 7112 27710 7168
rect 27766 7112 28262 7168
rect 28318 7112 28323 7168
rect 27705 7110 28323 7112
rect 27705 7107 27771 7110
rect 28257 7107 28323 7110
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 28441 6898 28507 6901
rect 28809 6898 28875 6901
rect 28441 6896 28875 6898
rect 28441 6840 28446 6896
rect 28502 6840 28814 6896
rect 28870 6840 28875 6896
rect 28441 6838 28875 6840
rect 28441 6835 28507 6838
rect 28809 6835 28875 6838
rect 27429 6762 27495 6765
rect 27981 6762 28047 6765
rect 28625 6762 28691 6765
rect 27429 6760 28691 6762
rect 27429 6704 27434 6760
rect 27490 6704 27986 6760
rect 28042 6704 28630 6760
rect 28686 6704 28691 6760
rect 27429 6702 28691 6704
rect 27429 6699 27495 6702
rect 27981 6699 28047 6702
rect 28625 6699 28691 6702
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 35590 6560 35906 6561
rect 35590 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35906 6560
rect 35590 6495 35906 6496
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 35590 5472 35906 5473
rect 35590 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35906 5472
rect 35590 5407 35906 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 35590 4384 35906 4385
rect 35590 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35906 4384
rect 35590 4319 35906 4320
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 35590 3296 35906 3297
rect 35590 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35906 3296
rect 35590 3231 35906 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 4870 2208 5186 2209
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 35590 2208 35906 2209
rect 35590 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35906 2208
rect 35590 2143 35906 2144
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 35596 37020 35660 37024
rect 35596 36964 35600 37020
rect 35600 36964 35656 37020
rect 35656 36964 35660 37020
rect 35596 36960 35660 36964
rect 35676 37020 35740 37024
rect 35676 36964 35680 37020
rect 35680 36964 35736 37020
rect 35736 36964 35740 37020
rect 35676 36960 35740 36964
rect 35756 37020 35820 37024
rect 35756 36964 35760 37020
rect 35760 36964 35816 37020
rect 35816 36964 35820 37020
rect 35756 36960 35820 36964
rect 35836 37020 35900 37024
rect 35836 36964 35840 37020
rect 35840 36964 35896 37020
rect 35896 36964 35900 37020
rect 35836 36960 35900 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 35596 35932 35660 35936
rect 35596 35876 35600 35932
rect 35600 35876 35656 35932
rect 35656 35876 35660 35932
rect 35596 35872 35660 35876
rect 35676 35932 35740 35936
rect 35676 35876 35680 35932
rect 35680 35876 35736 35932
rect 35736 35876 35740 35932
rect 35676 35872 35740 35876
rect 35756 35932 35820 35936
rect 35756 35876 35760 35932
rect 35760 35876 35816 35932
rect 35816 35876 35820 35932
rect 35756 35872 35820 35876
rect 35836 35932 35900 35936
rect 35836 35876 35840 35932
rect 35840 35876 35896 35932
rect 35896 35876 35900 35932
rect 35836 35872 35900 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 35596 34844 35660 34848
rect 35596 34788 35600 34844
rect 35600 34788 35656 34844
rect 35656 34788 35660 34844
rect 35596 34784 35660 34788
rect 35676 34844 35740 34848
rect 35676 34788 35680 34844
rect 35680 34788 35736 34844
rect 35736 34788 35740 34844
rect 35676 34784 35740 34788
rect 35756 34844 35820 34848
rect 35756 34788 35760 34844
rect 35760 34788 35816 34844
rect 35816 34788 35820 34844
rect 35756 34784 35820 34788
rect 35836 34844 35900 34848
rect 35836 34788 35840 34844
rect 35840 34788 35896 34844
rect 35896 34788 35900 34844
rect 35836 34784 35900 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 35596 33756 35660 33760
rect 35596 33700 35600 33756
rect 35600 33700 35656 33756
rect 35656 33700 35660 33756
rect 35596 33696 35660 33700
rect 35676 33756 35740 33760
rect 35676 33700 35680 33756
rect 35680 33700 35736 33756
rect 35736 33700 35740 33756
rect 35676 33696 35740 33700
rect 35756 33756 35820 33760
rect 35756 33700 35760 33756
rect 35760 33700 35816 33756
rect 35816 33700 35820 33756
rect 35756 33696 35820 33700
rect 35836 33756 35900 33760
rect 35836 33700 35840 33756
rect 35840 33700 35896 33756
rect 35896 33700 35900 33756
rect 35836 33696 35900 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 35596 32668 35660 32672
rect 35596 32612 35600 32668
rect 35600 32612 35656 32668
rect 35656 32612 35660 32668
rect 35596 32608 35660 32612
rect 35676 32668 35740 32672
rect 35676 32612 35680 32668
rect 35680 32612 35736 32668
rect 35736 32612 35740 32668
rect 35676 32608 35740 32612
rect 35756 32668 35820 32672
rect 35756 32612 35760 32668
rect 35760 32612 35816 32668
rect 35816 32612 35820 32668
rect 35756 32608 35820 32612
rect 35836 32668 35900 32672
rect 35836 32612 35840 32668
rect 35840 32612 35896 32668
rect 35896 32612 35900 32668
rect 35836 32608 35900 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 35596 31580 35660 31584
rect 35596 31524 35600 31580
rect 35600 31524 35656 31580
rect 35656 31524 35660 31580
rect 35596 31520 35660 31524
rect 35676 31580 35740 31584
rect 35676 31524 35680 31580
rect 35680 31524 35736 31580
rect 35736 31524 35740 31580
rect 35676 31520 35740 31524
rect 35756 31580 35820 31584
rect 35756 31524 35760 31580
rect 35760 31524 35816 31580
rect 35816 31524 35820 31580
rect 35756 31520 35820 31524
rect 35836 31580 35900 31584
rect 35836 31524 35840 31580
rect 35840 31524 35896 31580
rect 35896 31524 35900 31580
rect 35836 31520 35900 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 35596 30492 35660 30496
rect 35596 30436 35600 30492
rect 35600 30436 35656 30492
rect 35656 30436 35660 30492
rect 35596 30432 35660 30436
rect 35676 30492 35740 30496
rect 35676 30436 35680 30492
rect 35680 30436 35736 30492
rect 35736 30436 35740 30492
rect 35676 30432 35740 30436
rect 35756 30492 35820 30496
rect 35756 30436 35760 30492
rect 35760 30436 35816 30492
rect 35816 30436 35820 30492
rect 35756 30432 35820 30436
rect 35836 30492 35900 30496
rect 35836 30436 35840 30492
rect 35840 30436 35896 30492
rect 35896 30436 35900 30492
rect 35836 30432 35900 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 35596 29404 35660 29408
rect 35596 29348 35600 29404
rect 35600 29348 35656 29404
rect 35656 29348 35660 29404
rect 35596 29344 35660 29348
rect 35676 29404 35740 29408
rect 35676 29348 35680 29404
rect 35680 29348 35736 29404
rect 35736 29348 35740 29404
rect 35676 29344 35740 29348
rect 35756 29404 35820 29408
rect 35756 29348 35760 29404
rect 35760 29348 35816 29404
rect 35816 29348 35820 29404
rect 35756 29344 35820 29348
rect 35836 29404 35900 29408
rect 35836 29348 35840 29404
rect 35840 29348 35896 29404
rect 35896 29348 35900 29404
rect 35836 29344 35900 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 35596 28316 35660 28320
rect 35596 28260 35600 28316
rect 35600 28260 35656 28316
rect 35656 28260 35660 28316
rect 35596 28256 35660 28260
rect 35676 28316 35740 28320
rect 35676 28260 35680 28316
rect 35680 28260 35736 28316
rect 35736 28260 35740 28316
rect 35676 28256 35740 28260
rect 35756 28316 35820 28320
rect 35756 28260 35760 28316
rect 35760 28260 35816 28316
rect 35816 28260 35820 28316
rect 35756 28256 35820 28260
rect 35836 28316 35900 28320
rect 35836 28260 35840 28316
rect 35840 28260 35896 28316
rect 35896 28260 35900 28316
rect 35836 28256 35900 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 35596 27228 35660 27232
rect 35596 27172 35600 27228
rect 35600 27172 35656 27228
rect 35656 27172 35660 27228
rect 35596 27168 35660 27172
rect 35676 27228 35740 27232
rect 35676 27172 35680 27228
rect 35680 27172 35736 27228
rect 35736 27172 35740 27228
rect 35676 27168 35740 27172
rect 35756 27228 35820 27232
rect 35756 27172 35760 27228
rect 35760 27172 35816 27228
rect 35816 27172 35820 27228
rect 35756 27168 35820 27172
rect 35836 27228 35900 27232
rect 35836 27172 35840 27228
rect 35840 27172 35896 27228
rect 35896 27172 35900 27228
rect 35836 27168 35900 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 35596 26140 35660 26144
rect 35596 26084 35600 26140
rect 35600 26084 35656 26140
rect 35656 26084 35660 26140
rect 35596 26080 35660 26084
rect 35676 26140 35740 26144
rect 35676 26084 35680 26140
rect 35680 26084 35736 26140
rect 35736 26084 35740 26140
rect 35676 26080 35740 26084
rect 35756 26140 35820 26144
rect 35756 26084 35760 26140
rect 35760 26084 35816 26140
rect 35816 26084 35820 26140
rect 35756 26080 35820 26084
rect 35836 26140 35900 26144
rect 35836 26084 35840 26140
rect 35840 26084 35896 26140
rect 35896 26084 35900 26140
rect 35836 26080 35900 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 35596 25052 35660 25056
rect 35596 24996 35600 25052
rect 35600 24996 35656 25052
rect 35656 24996 35660 25052
rect 35596 24992 35660 24996
rect 35676 25052 35740 25056
rect 35676 24996 35680 25052
rect 35680 24996 35736 25052
rect 35736 24996 35740 25052
rect 35676 24992 35740 24996
rect 35756 25052 35820 25056
rect 35756 24996 35760 25052
rect 35760 24996 35816 25052
rect 35816 24996 35820 25052
rect 35756 24992 35820 24996
rect 35836 25052 35900 25056
rect 35836 24996 35840 25052
rect 35840 24996 35896 25052
rect 35896 24996 35900 25052
rect 35836 24992 35900 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 35596 23964 35660 23968
rect 35596 23908 35600 23964
rect 35600 23908 35656 23964
rect 35656 23908 35660 23964
rect 35596 23904 35660 23908
rect 35676 23964 35740 23968
rect 35676 23908 35680 23964
rect 35680 23908 35736 23964
rect 35736 23908 35740 23964
rect 35676 23904 35740 23908
rect 35756 23964 35820 23968
rect 35756 23908 35760 23964
rect 35760 23908 35816 23964
rect 35816 23908 35820 23964
rect 35756 23904 35820 23908
rect 35836 23964 35900 23968
rect 35836 23908 35840 23964
rect 35840 23908 35896 23964
rect 35896 23908 35900 23964
rect 35836 23904 35900 23908
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 35596 22876 35660 22880
rect 35596 22820 35600 22876
rect 35600 22820 35656 22876
rect 35656 22820 35660 22876
rect 35596 22816 35660 22820
rect 35676 22876 35740 22880
rect 35676 22820 35680 22876
rect 35680 22820 35736 22876
rect 35736 22820 35740 22876
rect 35676 22816 35740 22820
rect 35756 22876 35820 22880
rect 35756 22820 35760 22876
rect 35760 22820 35816 22876
rect 35816 22820 35820 22876
rect 35756 22816 35820 22820
rect 35836 22876 35900 22880
rect 35836 22820 35840 22876
rect 35840 22820 35896 22876
rect 35896 22820 35900 22876
rect 35836 22816 35900 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 35596 21788 35660 21792
rect 35596 21732 35600 21788
rect 35600 21732 35656 21788
rect 35656 21732 35660 21788
rect 35596 21728 35660 21732
rect 35676 21788 35740 21792
rect 35676 21732 35680 21788
rect 35680 21732 35736 21788
rect 35736 21732 35740 21788
rect 35676 21728 35740 21732
rect 35756 21788 35820 21792
rect 35756 21732 35760 21788
rect 35760 21732 35816 21788
rect 35816 21732 35820 21788
rect 35756 21728 35820 21732
rect 35836 21788 35900 21792
rect 35836 21732 35840 21788
rect 35840 21732 35896 21788
rect 35896 21732 35900 21788
rect 35836 21728 35900 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 34652 20980 34716 21044
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 35596 20700 35660 20704
rect 35596 20644 35600 20700
rect 35600 20644 35656 20700
rect 35656 20644 35660 20700
rect 35596 20640 35660 20644
rect 35676 20700 35740 20704
rect 35676 20644 35680 20700
rect 35680 20644 35736 20700
rect 35736 20644 35740 20700
rect 35676 20640 35740 20644
rect 35756 20700 35820 20704
rect 35756 20644 35760 20700
rect 35760 20644 35816 20700
rect 35816 20644 35820 20700
rect 35756 20640 35820 20644
rect 35836 20700 35900 20704
rect 35836 20644 35840 20700
rect 35840 20644 35896 20700
rect 35896 20644 35900 20700
rect 35836 20640 35900 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 35596 19612 35660 19616
rect 35596 19556 35600 19612
rect 35600 19556 35656 19612
rect 35656 19556 35660 19612
rect 35596 19552 35660 19556
rect 35676 19612 35740 19616
rect 35676 19556 35680 19612
rect 35680 19556 35736 19612
rect 35736 19556 35740 19612
rect 35676 19552 35740 19556
rect 35756 19612 35820 19616
rect 35756 19556 35760 19612
rect 35760 19556 35816 19612
rect 35816 19556 35820 19612
rect 35756 19552 35820 19556
rect 35836 19612 35900 19616
rect 35836 19556 35840 19612
rect 35840 19556 35896 19612
rect 35896 19556 35900 19612
rect 35836 19552 35900 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 35596 18524 35660 18528
rect 35596 18468 35600 18524
rect 35600 18468 35656 18524
rect 35656 18468 35660 18524
rect 35596 18464 35660 18468
rect 35676 18524 35740 18528
rect 35676 18468 35680 18524
rect 35680 18468 35736 18524
rect 35736 18468 35740 18524
rect 35676 18464 35740 18468
rect 35756 18524 35820 18528
rect 35756 18468 35760 18524
rect 35760 18468 35816 18524
rect 35816 18468 35820 18524
rect 35756 18464 35820 18468
rect 35836 18524 35900 18528
rect 35836 18468 35840 18524
rect 35840 18468 35896 18524
rect 35896 18468 35900 18524
rect 35836 18464 35900 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 35596 17436 35660 17440
rect 35596 17380 35600 17436
rect 35600 17380 35656 17436
rect 35656 17380 35660 17436
rect 35596 17376 35660 17380
rect 35676 17436 35740 17440
rect 35676 17380 35680 17436
rect 35680 17380 35736 17436
rect 35736 17380 35740 17436
rect 35676 17376 35740 17380
rect 35756 17436 35820 17440
rect 35756 17380 35760 17436
rect 35760 17380 35816 17436
rect 35816 17380 35820 17436
rect 35756 17376 35820 17380
rect 35836 17436 35900 17440
rect 35836 17380 35840 17436
rect 35840 17380 35896 17436
rect 35896 17380 35900 17436
rect 35836 17376 35900 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 35596 16348 35660 16352
rect 35596 16292 35600 16348
rect 35600 16292 35656 16348
rect 35656 16292 35660 16348
rect 35596 16288 35660 16292
rect 35676 16348 35740 16352
rect 35676 16292 35680 16348
rect 35680 16292 35736 16348
rect 35736 16292 35740 16348
rect 35676 16288 35740 16292
rect 35756 16348 35820 16352
rect 35756 16292 35760 16348
rect 35760 16292 35816 16348
rect 35816 16292 35820 16348
rect 35756 16288 35820 16292
rect 35836 16348 35900 16352
rect 35836 16292 35840 16348
rect 35840 16292 35896 16348
rect 35896 16292 35900 16348
rect 35836 16288 35900 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 35596 15260 35660 15264
rect 35596 15204 35600 15260
rect 35600 15204 35656 15260
rect 35656 15204 35660 15260
rect 35596 15200 35660 15204
rect 35676 15260 35740 15264
rect 35676 15204 35680 15260
rect 35680 15204 35736 15260
rect 35736 15204 35740 15260
rect 35676 15200 35740 15204
rect 35756 15260 35820 15264
rect 35756 15204 35760 15260
rect 35760 15204 35816 15260
rect 35816 15204 35820 15260
rect 35756 15200 35820 15204
rect 35836 15260 35900 15264
rect 35836 15204 35840 15260
rect 35840 15204 35896 15260
rect 35896 15204 35900 15260
rect 35836 15200 35900 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 35596 14172 35660 14176
rect 35596 14116 35600 14172
rect 35600 14116 35656 14172
rect 35656 14116 35660 14172
rect 35596 14112 35660 14116
rect 35676 14172 35740 14176
rect 35676 14116 35680 14172
rect 35680 14116 35736 14172
rect 35736 14116 35740 14172
rect 35676 14112 35740 14116
rect 35756 14172 35820 14176
rect 35756 14116 35760 14172
rect 35760 14116 35816 14172
rect 35816 14116 35820 14172
rect 35756 14112 35820 14116
rect 35836 14172 35900 14176
rect 35836 14116 35840 14172
rect 35840 14116 35896 14172
rect 35896 14116 35900 14172
rect 35836 14112 35900 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 35596 13084 35660 13088
rect 35596 13028 35600 13084
rect 35600 13028 35656 13084
rect 35656 13028 35660 13084
rect 35596 13024 35660 13028
rect 35676 13084 35740 13088
rect 35676 13028 35680 13084
rect 35680 13028 35736 13084
rect 35736 13028 35740 13084
rect 35676 13024 35740 13028
rect 35756 13084 35820 13088
rect 35756 13028 35760 13084
rect 35760 13028 35816 13084
rect 35816 13028 35820 13084
rect 35756 13024 35820 13028
rect 35836 13084 35900 13088
rect 35836 13028 35840 13084
rect 35840 13028 35896 13084
rect 35896 13028 35900 13084
rect 35836 13024 35900 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 35596 11996 35660 12000
rect 35596 11940 35600 11996
rect 35600 11940 35656 11996
rect 35656 11940 35660 11996
rect 35596 11936 35660 11940
rect 35676 11996 35740 12000
rect 35676 11940 35680 11996
rect 35680 11940 35736 11996
rect 35736 11940 35740 11996
rect 35676 11936 35740 11940
rect 35756 11996 35820 12000
rect 35756 11940 35760 11996
rect 35760 11940 35816 11996
rect 35816 11940 35820 11996
rect 35756 11936 35820 11940
rect 35836 11996 35900 12000
rect 35836 11940 35840 11996
rect 35840 11940 35896 11996
rect 35896 11940 35900 11996
rect 35836 11936 35900 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 34652 10916 34716 10980
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 35596 10908 35660 10912
rect 35596 10852 35600 10908
rect 35600 10852 35656 10908
rect 35656 10852 35660 10908
rect 35596 10848 35660 10852
rect 35676 10908 35740 10912
rect 35676 10852 35680 10908
rect 35680 10852 35736 10908
rect 35736 10852 35740 10908
rect 35676 10848 35740 10852
rect 35756 10908 35820 10912
rect 35756 10852 35760 10908
rect 35760 10852 35816 10908
rect 35816 10852 35820 10908
rect 35756 10848 35820 10852
rect 35836 10908 35900 10912
rect 35836 10852 35840 10908
rect 35840 10852 35896 10908
rect 35896 10852 35900 10908
rect 35836 10848 35900 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 35596 9820 35660 9824
rect 35596 9764 35600 9820
rect 35600 9764 35656 9820
rect 35656 9764 35660 9820
rect 35596 9760 35660 9764
rect 35676 9820 35740 9824
rect 35676 9764 35680 9820
rect 35680 9764 35736 9820
rect 35736 9764 35740 9820
rect 35676 9760 35740 9764
rect 35756 9820 35820 9824
rect 35756 9764 35760 9820
rect 35760 9764 35816 9820
rect 35816 9764 35820 9820
rect 35756 9760 35820 9764
rect 35836 9820 35900 9824
rect 35836 9764 35840 9820
rect 35840 9764 35896 9820
rect 35896 9764 35900 9820
rect 35836 9760 35900 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 35596 8732 35660 8736
rect 35596 8676 35600 8732
rect 35600 8676 35656 8732
rect 35656 8676 35660 8732
rect 35596 8672 35660 8676
rect 35676 8732 35740 8736
rect 35676 8676 35680 8732
rect 35680 8676 35736 8732
rect 35736 8676 35740 8732
rect 35676 8672 35740 8676
rect 35756 8732 35820 8736
rect 35756 8676 35760 8732
rect 35760 8676 35816 8732
rect 35816 8676 35820 8732
rect 35756 8672 35820 8676
rect 35836 8732 35900 8736
rect 35836 8676 35840 8732
rect 35840 8676 35896 8732
rect 35896 8676 35900 8732
rect 35836 8672 35900 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 35596 7644 35660 7648
rect 35596 7588 35600 7644
rect 35600 7588 35656 7644
rect 35656 7588 35660 7644
rect 35596 7584 35660 7588
rect 35676 7644 35740 7648
rect 35676 7588 35680 7644
rect 35680 7588 35736 7644
rect 35736 7588 35740 7644
rect 35676 7584 35740 7588
rect 35756 7644 35820 7648
rect 35756 7588 35760 7644
rect 35760 7588 35816 7644
rect 35816 7588 35820 7644
rect 35756 7584 35820 7588
rect 35836 7644 35900 7648
rect 35836 7588 35840 7644
rect 35840 7588 35896 7644
rect 35896 7588 35900 7644
rect 35836 7584 35900 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 35596 6556 35660 6560
rect 35596 6500 35600 6556
rect 35600 6500 35656 6556
rect 35656 6500 35660 6556
rect 35596 6496 35660 6500
rect 35676 6556 35740 6560
rect 35676 6500 35680 6556
rect 35680 6500 35736 6556
rect 35736 6500 35740 6556
rect 35676 6496 35740 6500
rect 35756 6556 35820 6560
rect 35756 6500 35760 6556
rect 35760 6500 35816 6556
rect 35816 6500 35820 6556
rect 35756 6496 35820 6500
rect 35836 6556 35900 6560
rect 35836 6500 35840 6556
rect 35840 6500 35896 6556
rect 35896 6500 35900 6556
rect 35836 6496 35900 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 35596 5468 35660 5472
rect 35596 5412 35600 5468
rect 35600 5412 35656 5468
rect 35656 5412 35660 5468
rect 35596 5408 35660 5412
rect 35676 5468 35740 5472
rect 35676 5412 35680 5468
rect 35680 5412 35736 5468
rect 35736 5412 35740 5468
rect 35676 5408 35740 5412
rect 35756 5468 35820 5472
rect 35756 5412 35760 5468
rect 35760 5412 35816 5468
rect 35816 5412 35820 5468
rect 35756 5408 35820 5412
rect 35836 5468 35900 5472
rect 35836 5412 35840 5468
rect 35840 5412 35896 5468
rect 35896 5412 35900 5468
rect 35836 5408 35900 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 35596 4380 35660 4384
rect 35596 4324 35600 4380
rect 35600 4324 35656 4380
rect 35656 4324 35660 4380
rect 35596 4320 35660 4324
rect 35676 4380 35740 4384
rect 35676 4324 35680 4380
rect 35680 4324 35736 4380
rect 35736 4324 35740 4380
rect 35676 4320 35740 4324
rect 35756 4380 35820 4384
rect 35756 4324 35760 4380
rect 35760 4324 35816 4380
rect 35816 4324 35820 4380
rect 35756 4320 35820 4324
rect 35836 4380 35900 4384
rect 35836 4324 35840 4380
rect 35840 4324 35896 4380
rect 35896 4324 35900 4380
rect 35836 4320 35900 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 35596 3292 35660 3296
rect 35596 3236 35600 3292
rect 35600 3236 35656 3292
rect 35656 3236 35660 3292
rect 35596 3232 35660 3236
rect 35676 3292 35740 3296
rect 35676 3236 35680 3292
rect 35680 3236 35736 3292
rect 35736 3236 35740 3292
rect 35676 3232 35740 3236
rect 35756 3292 35820 3296
rect 35756 3236 35760 3292
rect 35760 3236 35816 3292
rect 35816 3236 35820 3292
rect 35756 3232 35820 3236
rect 35836 3292 35900 3296
rect 35836 3236 35840 3292
rect 35840 3236 35896 3292
rect 35896 3236 35900 3292
rect 35836 3232 35900 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
rect 35596 2204 35660 2208
rect 35596 2148 35600 2204
rect 35600 2148 35656 2204
rect 35656 2148 35660 2204
rect 35596 2144 35660 2148
rect 35676 2204 35740 2208
rect 35676 2148 35680 2204
rect 35680 2148 35736 2204
rect 35736 2148 35740 2204
rect 35676 2144 35740 2148
rect 35756 2204 35820 2208
rect 35756 2148 35760 2204
rect 35760 2148 35816 2204
rect 35816 2148 35820 2204
rect 35756 2144 35820 2148
rect 35836 2204 35900 2208
rect 35836 2148 35840 2204
rect 35840 2148 35896 2204
rect 35896 2148 35900 2204
rect 35836 2144 35900 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36260 4528 36416
rect 4208 36024 4250 36260
rect 4486 36024 4528 36260
rect 4208 35392 4528 36024
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5624 4528 5952
rect 4208 5388 4250 5624
rect 4486 5388 4528 5624
rect 4208 4928 4528 5388
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 37024 5188 37584
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 4868 36920 5188 36960
rect 4868 36684 4910 36920
rect 5146 36684 5188 36920
rect 4868 35936 5188 36684
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36260 35248 36416
rect 34928 36024 34970 36260
rect 35206 36024 35248 36260
rect 34928 35392 35248 36024
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34651 21044 34717 21045
rect 34651 20980 34652 21044
rect 34716 20980 34717 21044
rect 34651 20979 34717 20980
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 34654 10981 34714 20979
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34651 10980 34717 10981
rect 34651 10916 34652 10980
rect 34716 10916 34717 10980
rect 34651 10915 34717 10916
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 6284 5188 6496
rect 4868 6048 4910 6284
rect 5146 6048 5188 6284
rect 4868 5472 5188 6048
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5624 35248 5952
rect 34928 5388 34970 5624
rect 35206 5388 35248 5624
rect 34928 4928 35248 5388
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 35588 37024 35908 37584
rect 35588 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35908 37024
rect 35588 36920 35908 36960
rect 35588 36684 35630 36920
rect 35866 36684 35908 36920
rect 35588 35936 35908 36684
rect 35588 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35908 35936
rect 35588 34848 35908 35872
rect 35588 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35908 34848
rect 35588 33760 35908 34784
rect 35588 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35908 33760
rect 35588 32672 35908 33696
rect 35588 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35908 32672
rect 35588 31584 35908 32608
rect 35588 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35908 31584
rect 35588 30496 35908 31520
rect 35588 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35908 30496
rect 35588 29408 35908 30432
rect 35588 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35908 29408
rect 35588 28320 35908 29344
rect 35588 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35908 28320
rect 35588 27232 35908 28256
rect 35588 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35908 27232
rect 35588 26144 35908 27168
rect 35588 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35908 26144
rect 35588 25056 35908 26080
rect 35588 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35908 25056
rect 35588 23968 35908 24992
rect 35588 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35908 23968
rect 35588 22880 35908 23904
rect 35588 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35908 22880
rect 35588 21792 35908 22816
rect 35588 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35908 21792
rect 35588 20704 35908 21728
rect 35588 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35908 20704
rect 35588 19616 35908 20640
rect 35588 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35908 19616
rect 35588 18528 35908 19552
rect 35588 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35908 18528
rect 35588 17440 35908 18464
rect 35588 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35908 17440
rect 35588 16352 35908 17376
rect 35588 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35908 16352
rect 35588 15264 35908 16288
rect 35588 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35908 15264
rect 35588 14176 35908 15200
rect 35588 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35908 14176
rect 35588 13088 35908 14112
rect 35588 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35908 13088
rect 35588 12000 35908 13024
rect 35588 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35908 12000
rect 35588 10912 35908 11936
rect 35588 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35908 10912
rect 35588 9824 35908 10848
rect 35588 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35908 9824
rect 35588 8736 35908 9760
rect 35588 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35908 8736
rect 35588 7648 35908 8672
rect 35588 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35908 7648
rect 35588 6560 35908 7584
rect 35588 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35908 6560
rect 35588 6284 35908 6496
rect 35588 6048 35630 6284
rect 35866 6048 35908 6284
rect 35588 5472 35908 6048
rect 35588 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35908 5472
rect 35588 4384 35908 5408
rect 35588 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35908 4384
rect 35588 3296 35908 4320
rect 35588 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35908 3296
rect 35588 2208 35908 3232
rect 35588 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35908 2208
rect 35588 2128 35908 2144
<< via4 >>
rect 4250 36024 4486 36260
rect 4250 5388 4486 5624
rect 4910 36684 5146 36920
rect 34970 36024 35206 36260
rect 4910 6048 5146 6284
rect 34970 5388 35206 5624
rect 35630 36684 35866 36920
rect 35630 6048 35866 6284
<< metal5 >>
rect 1056 36920 38872 36962
rect 1056 36684 4910 36920
rect 5146 36684 35630 36920
rect 35866 36684 38872 36920
rect 1056 36642 38872 36684
rect 1056 36260 38872 36302
rect 1056 36024 4250 36260
rect 4486 36024 34970 36260
rect 35206 36024 38872 36260
rect 1056 35982 38872 36024
rect 1056 6284 38872 6326
rect 1056 6048 4910 6284
rect 5146 6048 35630 6284
rect 35866 6048 38872 6284
rect 1056 6006 38872 6048
rect 1056 5624 38872 5666
rect 1056 5388 4250 5624
rect 4486 5388 34970 5624
rect 35206 5388 38872 5624
rect 1056 5346 38872 5388
use sky130_fd_sc_hd__xnor2_1  _112_
timestamp 0
transform 1 0 23460 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _113_
timestamp 0
transform 1 0 23184 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _114_
timestamp 0
transform 1 0 24380 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _115_
timestamp 0
transform 1 0 20240 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _116_
timestamp 0
transform 1 0 19228 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _117_
timestamp 0
transform 1 0 21804 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _118_
timestamp 0
transform 1 0 24840 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _119_
timestamp 0
transform 1 0 29624 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor3_2  _120_
timestamp 0
transform 1 0 26772 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _121_
timestamp 0
transform -1 0 28428 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _122_
timestamp 0
transform 1 0 25300 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 0
transform 1 0 25484 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _124_
timestamp 0
transform -1 0 27784 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  _125_
timestamp 0
transform -1 0 25668 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__or2_1  _126_
timestamp 0
transform 1 0 23828 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__mux4_1  _127_
timestamp 0
transform 1 0 21804 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__or2b_1  _128_
timestamp 0
transform 1 0 24472 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _129_
timestamp 0
transform -1 0 26864 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _130_
timestamp 0
transform -1 0 27416 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _131_
timestamp 0
transform 1 0 25208 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _132_
timestamp 0
transform 1 0 25944 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _133_
timestamp 0
transform 1 0 25392 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _134_
timestamp 0
transform -1 0 27600 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _135_
timestamp 0
transform -1 0 27968 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _136_
timestamp 0
transform 1 0 28520 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _137_
timestamp 0
transform 1 0 26956 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _138_
timestamp 0
transform 1 0 23552 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _139_
timestamp 0
transform 1 0 22908 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _140_
timestamp 0
transform -1 0 30084 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _141_
timestamp 0
transform -1 0 28980 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _142_
timestamp 0
transform 1 0 25852 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _143_
timestamp 0
transform -1 0 25944 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _144_
timestamp 0
transform -1 0 25024 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _145_
timestamp 0
transform -1 0 29164 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _146_
timestamp 0
transform 1 0 26036 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _147_
timestamp 0
transform -1 0 26864 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _148_
timestamp 0
transform 1 0 27968 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _149_
timestamp 0
transform 1 0 26312 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and4_1  _150_
timestamp 0
transform 1 0 26496 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and4b_1  _151_
timestamp 0
transform 1 0 26956 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _152_
timestamp 0
transform 1 0 27876 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _153_
timestamp 0
transform -1 0 27876 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _154_
timestamp 0
transform -1 0 26036 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _155_
timestamp 0
transform -1 0 26864 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _156_
timestamp 0
transform -1 0 26036 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _157_
timestamp 0
transform 1 0 24840 0 1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 0
transform 1 0 24564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _159_
timestamp 0
transform 1 0 26956 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _160_
timestamp 0
transform -1 0 26864 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _161_
timestamp 0
transform 1 0 25944 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _162_
timestamp 0
transform 1 0 26404 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _163_
timestamp 0
transform -1 0 26864 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _164_
timestamp 0
transform 1 0 25668 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _165_
timestamp 0
transform 1 0 28428 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _166_
timestamp 0
transform -1 0 27600 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _167_
timestamp 0
transform -1 0 28520 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _168_
timestamp 0
transform 1 0 28888 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _169_
timestamp 0
transform 1 0 27876 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _170_
timestamp 0
transform -1 0 28520 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_1  _171_
timestamp 0
transform 1 0 29532 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _172_
timestamp 0
transform -1 0 30636 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _173_
timestamp 0
transform 1 0 28336 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _174_
timestamp 0
transform 1 0 29532 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _175_
timestamp 0
transform 1 0 27600 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _176_
timestamp 0
transform -1 0 28060 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_1  _177_
timestamp 0
transform 1 0 25944 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _178_
timestamp 0
transform 1 0 27692 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _179_
timestamp 0
transform 1 0 29532 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _180_
timestamp 0
transform 1 0 26956 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _181_
timestamp 0
transform -1 0 27692 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _182_
timestamp 0
transform -1 0 28520 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _183_
timestamp 0
transform -1 0 22540 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _184_
timestamp 0
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _185_
timestamp 0
transform -1 0 25116 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _186_
timestamp 0
transform -1 0 24196 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _187_
timestamp 0
transform 1 0 20792 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _188_
timestamp 0
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _189_
timestamp 0
transform -1 0 24840 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _190_
timestamp 0
transform 1 0 22448 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _191_
timestamp 0
transform -1 0 24564 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _192_
timestamp 0
transform -1 0 23552 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _193_
timestamp 0
transform -1 0 21712 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _194_
timestamp 0
transform 1 0 20516 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _195_
timestamp 0
transform -1 0 24104 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _196_
timestamp 0
transform 1 0 22632 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _197_
timestamp 0
transform -1 0 25576 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _198_
timestamp 0
transform -1 0 25392 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _199_
timestamp 0
transform 1 0 25576 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _200_
timestamp 0
transform 1 0 21804 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _201_
timestamp 0
transform 1 0 21252 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _202_
timestamp 0
transform 1 0 22632 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _203_
timestamp 0
transform -1 0 23920 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _204_
timestamp 0
transform 1 0 22816 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _205_
timestamp 0
transform -1 0 25852 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o2111a_1  _206_
timestamp 0
transform 1 0 24380 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_1  _207_
timestamp 0
transform 1 0 23736 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _208_
timestamp 0
transform 1 0 23460 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _209_
timestamp 0
transform 1 0 23184 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _210_
timestamp 0
transform 1 0 23276 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _211_
timestamp 0
transform 1 0 22908 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _212_
timestamp 0
transform 1 0 19228 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _213_
timestamp 0
transform 1 0 18768 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _214_
timestamp 0
transform 1 0 18308 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _215_
timestamp 0
transform -1 0 18308 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _216_
timestamp 0
transform 1 0 21528 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _217_
timestamp 0
transform 1 0 21252 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _218_
timestamp 0
transform 1 0 19412 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _219_
timestamp 0
transform -1 0 19412 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _220_
timestamp 0
transform 1 0 21804 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _221_
timestamp 0
transform 1 0 20516 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _222_
timestamp 0
transform 1 0 21620 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _223_
timestamp 0
transform 1 0 21160 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _224_
timestamp 0
transform 1 0 24840 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _225_
timestamp 0
transform 1 0 24840 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _226_
timestamp 0
transform -1 0 28244 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _227_
timestamp 0
transform 1 0 27416 0 -1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _228_
timestamp 0
transform 1 0 27784 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _229_
timestamp 0
transform 1 0 27508 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _230_
timestamp 0
transform 1 0 23736 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _231_
timestamp 0
transform 1 0 26220 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _232_
timestamp 0
transform 1 0 24380 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _233_
timestamp 0
transform -1 0 29532 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _234_
timestamp 0
transform 1 0 28520 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _235_
timestamp 0
transform -1 0 29992 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _236_
timestamp 0
transform 1 0 24104 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _237_
timestamp 0
transform -1 0 26220 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _238_
timestamp 0
transform 1 0 27416 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _239_
timestamp 0
transform 1 0 21160 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _240_
timestamp 0
transform -1 0 24656 0 -1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _241_
timestamp 0
transform 1 0 19872 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _242_
timestamp 0
transform 1 0 21896 0 -1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _243_
timestamp 0
transform -1 0 24012 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _244_
timestamp 0
transform 1 0 20148 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _245_
timestamp 0
transform 1 0 21804 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _246_
timestamp 0
transform 1 0 20700 0 1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _247_
timestamp 0
transform 1 0 21804 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _248_
timestamp 0
transform 1 0 23000 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _249_
timestamp 0
transform 1 0 22908 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _250_
timestamp 0
transform 1 0 22448 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _251_
timestamp 0
transform 1 0 18584 0 -1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _252_
timestamp 0
transform 1 0 18676 0 -1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _253_
timestamp 0
transform 1 0 20884 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _254_
timestamp 0
transform 1 0 19228 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _255_
timestamp 0
transform 1 0 19872 0 -1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _256_
timestamp 0
transform 1 0 20608 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 0
transform -1 0 26312 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 0
transform -1 0 22632 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 0
transform -1 0 22632 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 0
transform 1 0 26036 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 0
transform 1 0 26036 0 1 9792
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_4  fanout13
timestamp 0
transform -1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout14
timestamp 0
transform 1 0 21988 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  fanout15
timestamp 0
transform 1 0 25668 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  fanout16
timestamp 0
transform 1 0 25944 0 -1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_7
timestamp 0
transform 1 0 1748 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_19
timestamp 0
transform 1 0 2852 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 0
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 0
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_41
timestamp 0
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53
timestamp 0
transform 1 0 5980 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 0
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_69
timestamp 0
transform 1 0 7452 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81
timestamp 0
transform 1 0 8556 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 0
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_97
timestamp 0
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 0
transform 1 0 11132 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_113
timestamp 0
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_119
timestamp 0
transform 1 0 12052 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_131
timestamp 0
transform 1 0 13156 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 0
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_141
timestamp 0
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_153
timestamp 0
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 0
transform 1 0 16284 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 0
transform 1 0 16652 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_181
timestamp 0
transform 1 0 17756 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 0
transform 1 0 18860 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_197
timestamp 0
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_209
timestamp 0
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 0
transform 1 0 21436 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 0
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_237
timestamp 0
transform 1 0 22908 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_245
timestamp 0
transform 1 0 23644 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_251
timestamp 0
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 0
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 0
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 0
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 0
transform 1 0 26956 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 0
transform 1 0 28060 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 0
transform 1 0 29164 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 0
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 0
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 0
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_337
timestamp 0
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_349
timestamp 0
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 0
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_365
timestamp 0
transform 1 0 34684 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_373
timestamp 0
transform 1 0 35420 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_378
timestamp 0
transform 1 0 35880 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_390
timestamp 0
transform 1 0 36984 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_393
timestamp 0
transform 1 0 37260 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_405
timestamp 0
transform 1 0 38364 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 0
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 0
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 0
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 0
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 0
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 0
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 0
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 0
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 0
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 0
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 0
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 0
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 0
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 0
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 0
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 0
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 0
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 0
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 0
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 0
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 0
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 0
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 0
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 0
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 0
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 0
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 0
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 0
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 0
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 0
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 0
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 0
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 0
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 0
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 0
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 0
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 0
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 0
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_361
timestamp 0
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_373
timestamp 0
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_385
timestamp 0
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 0
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_393
timestamp 0
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_405
timestamp 0
transform 1 0 38364 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 0
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 0
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 0
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 0
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 0
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 0
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 0
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 0
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 0
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 0
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 0
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 0
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 0
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 0
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 0
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 0
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 0
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 0
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 0
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 0
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 0
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 0
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 0
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 0
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 0
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 0
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 0
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 0
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 0
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 0
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 0
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 0
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 0
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 0
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 0
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 0
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 0
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 0
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 0
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 0
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 0
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 0
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_401
timestamp 0
transform 1 0 37996 0 1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 0
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 0
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 0
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 0
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 0
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 0
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 0
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 0
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 0
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 0
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 0
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 0
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 0
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 0
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 0
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 0
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 0
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 0
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 0
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 0
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 0
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 0
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 0
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 0
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 0
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 0
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 0
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 0
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 0
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 0
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 0
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 0
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 0
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 0
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 0
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 0
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 0
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 0
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 0
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 0
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 0
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 0
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 0
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_405
timestamp 0
transform 1 0 38364 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 0
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 0
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 0
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 0
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 0
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 0
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 0
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 0
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 0
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 0
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 0
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 0
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 0
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 0
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 0
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 0
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 0
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 0
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 0
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 0
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 0
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 0
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 0
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 0
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 0
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 0
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 0
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 0
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 0
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_277
timestamp 0
transform 1 0 26588 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_287
timestamp 0
transform 1 0 27508 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_299
timestamp 0
transform 1 0 28612 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 0
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 0
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 0
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 0
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 0
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 0
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 0
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 0
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 0
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 0
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_401
timestamp 0
transform 1 0 37996 0 1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 0
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 0
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 0
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 0
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 0
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 0
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 0
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 0
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 0
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 0
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 0
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 0
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 0
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 0
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 0
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 0
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 0
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 0
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 0
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 0
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 0
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 0
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 0
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 0
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_225
timestamp 0
transform 1 0 21804 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_231
timestamp 0
transform 1 0 22356 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_235
timestamp 0
transform 1 0 22724 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_247
timestamp 0
transform 1 0 23828 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_259
timestamp 0
transform 1 0 24932 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_267
timestamp 0
transform 1 0 25668 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_278
timestamp 0
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_281
timestamp 0
transform 1 0 26956 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_291
timestamp 0
transform 1 0 27876 0 -1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_300
timestamp 0
transform 1 0 28704 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_312
timestamp 0
transform 1 0 29808 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_324
timestamp 0
transform 1 0 30912 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 0
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 0
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 0
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 0
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 0
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 0
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 0
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_405
timestamp 0
transform 1 0 38364 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 0
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 0
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 0
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 0
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 0
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 0
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 0
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 0
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 0
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 0
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 0
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 0
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 0
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 0
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 0
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 0
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 0
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 0
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 0
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 0
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 0
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 0
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 0
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_221
timestamp 0
transform 1 0 21436 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_249
timestamp 0
transform 1 0 24012 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_293
timestamp 0
transform 1 0 28060 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_306
timestamp 0
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 0
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 0
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 0
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 0
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 0
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 0
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 0
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 0
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 0
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_401
timestamp 0
transform 1 0 37996 0 1 5440
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 0
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 0
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 0
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 0
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 0
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 0
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 0
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 0
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 0
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 0
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 0
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 0
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 0
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 0
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 0
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 0
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 0
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 0
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 0
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 0
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_193
timestamp 0
transform 1 0 18860 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_201
timestamp 0
transform 1 0 19596 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_225
timestamp 0
transform 1 0 21804 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_309
timestamp 0
transform 1 0 29532 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_321
timestamp 0
transform 1 0 30636 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_333
timestamp 0
transform 1 0 31740 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 0
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 0
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 0
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 0
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 0
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 0
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 0
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_405
timestamp 0
transform 1 0 38364 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 0
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 0
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 0
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 0
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 0
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 0
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 0
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 0
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 0
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 0
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 0
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 0
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 0
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 0
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 0
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 0
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 0
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 0
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 0
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 0
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 0
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_197
timestamp 0
transform 1 0 19228 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_205
timestamp 0
transform 1 0 19964 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_288
timestamp 0
transform 1 0 27600 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_304
timestamp 0
transform 1 0 29072 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_315
timestamp 0
transform 1 0 30084 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_327
timestamp 0
transform 1 0 31188 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_339
timestamp 0
transform 1 0 32292 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_351
timestamp 0
transform 1 0 33396 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 0
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 0
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 0
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 0
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_401
timestamp 0
transform 1 0 37996 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 0
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 0
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 0
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 0
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 0
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 0
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 0
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 0
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 0
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 0
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 0
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 0
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 0
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 0
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 0
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 0
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 0
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 0
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 0
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 0
transform 1 0 17756 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 0
transform 1 0 18860 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_205
timestamp 0
transform 1 0 19964 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_258
timestamp 0
transform 1 0 24840 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_270
timestamp 0
transform 1 0 25944 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_318
timestamp 0
transform 1 0 30360 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_330
timestamp 0
transform 1 0 31464 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 0
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 0
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 0
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 0
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 0
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 0
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 0
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_405
timestamp 0
transform 1 0 38364 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 0
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 0
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 0
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 0
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 0
transform 1 0 4876 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 0
transform 1 0 5980 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 0
transform 1 0 7084 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 0
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 0
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 0
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 0
transform 1 0 10028 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 0
transform 1 0 11132 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 0
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 0
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 0
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 0
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 0
transform 1 0 15180 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 0
transform 1 0 16284 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 0
transform 1 0 17388 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 0
transform 1 0 18492 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 0
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 0
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_209
timestamp 0
transform 1 0 20332 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_213
timestamp 0
transform 1 0 20700 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 0
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 0
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_265
timestamp 0
transform 1 0 25484 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_304
timestamp 0
transform 1 0 29072 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_325
timestamp 0
transform 1 0 31004 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_337
timestamp 0
transform 1 0 32108 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_349
timestamp 0
transform 1 0 33212 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_361
timestamp 0
transform 1 0 34316 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 0
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 0
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 0
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_401
timestamp 0
transform 1 0 37996 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 0
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 0
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 0
transform 1 0 3588 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 0
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 0
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 0
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 0
transform 1 0 6348 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 0
transform 1 0 7452 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 0
transform 1 0 8556 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 0
transform 1 0 9660 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 0
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 0
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 0
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 0
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 0
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 0
transform 1 0 14812 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 0
transform 1 0 15916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 0
transform 1 0 16468 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_169
timestamp 0
transform 1 0 16652 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_181
timestamp 0
transform 1 0 17756 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_193
timestamp 0
transform 1 0 18860 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 0
transform 1 0 19964 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_217
timestamp 0
transform 1 0 21068 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_278
timestamp 0
transform 1 0 26680 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_293
timestamp 0
transform 1 0 28060 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_321
timestamp 0
transform 1 0 30636 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_333
timestamp 0
transform 1 0 31740 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 0
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 0
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_361
timestamp 0
transform 1 0 34316 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_373
timestamp 0
transform 1 0 35420 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_385
timestamp 0
transform 1 0 36524 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 0
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_393
timestamp 0
transform 1 0 37260 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_401
timestamp 0
transform 1 0 37996 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 0
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 0
transform 1 0 2484 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 0
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 0
transform 1 0 3772 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_41
timestamp 0
transform 1 0 4876 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_53
timestamp 0
transform 1 0 5980 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_65
timestamp 0
transform 1 0 7084 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_77
timestamp 0
transform 1 0 8188 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_83
timestamp 0
transform 1 0 8740 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_85
timestamp 0
transform 1 0 8924 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_97
timestamp 0
transform 1 0 10028 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_109
timestamp 0
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_121
timestamp 0
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_133
timestamp 0
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 0
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_141
timestamp 0
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_153
timestamp 0
transform 1 0 15180 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_165
timestamp 0
transform 1 0 16284 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_177
timestamp 0
transform 1 0 17388 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_189
timestamp 0
transform 1 0 18492 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_195
timestamp 0
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 0
transform 1 0 19228 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_209
timestamp 0
transform 1 0 20332 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_217
timestamp 0
transform 1 0 21068 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_238
timestamp 0
transform 1 0 23000 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 0
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_303
timestamp 0
transform 1 0 28980 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 0
transform 1 0 29348 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_315
timestamp 0
transform 1 0 30084 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_327
timestamp 0
transform 1 0 31188 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_339
timestamp 0
transform 1 0 32292 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_351
timestamp 0
transform 1 0 33396 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 0
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 0
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 0
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_389
timestamp 0
transform 1 0 36892 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_401
timestamp 0
transform 1 0 37996 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 0
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 0
transform 1 0 2484 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_27
timestamp 0
transform 1 0 3588 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_39
timestamp 0
transform 1 0 4692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 0
transform 1 0 5796 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 0
transform 1 0 6164 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_57
timestamp 0
transform 1 0 6348 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_69
timestamp 0
transform 1 0 7452 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_81
timestamp 0
transform 1 0 8556 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_93
timestamp 0
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_105
timestamp 0
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 0
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 0
transform 1 0 11500 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 0
transform 1 0 12604 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 0
transform 1 0 13708 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_149
timestamp 0
transform 1 0 14812 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_161
timestamp 0
transform 1 0 15916 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_167
timestamp 0
transform 1 0 16468 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_169
timestamp 0
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_181
timestamp 0
transform 1 0 17756 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_193
timestamp 0
transform 1 0 18860 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_205
timestamp 0
transform 1 0 19964 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_217
timestamp 0
transform 1 0 21068 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 0
transform 1 0 21620 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_225
timestamp 0
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_233
timestamp 0
transform 1 0 22540 0 -1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_306
timestamp 0
transform 1 0 29256 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_318
timestamp 0
transform 1 0 30360 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_330
timestamp 0
transform 1 0 31464 0 -1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_337
timestamp 0
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_349
timestamp 0
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_361
timestamp 0
transform 1 0 34316 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_373
timestamp 0
transform 1 0 35420 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_385
timestamp 0
transform 1 0 36524 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_391
timestamp 0
transform 1 0 37076 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_393
timestamp 0
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_405
timestamp 0
transform 1 0 38364 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 0
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_15
timestamp 0
transform 1 0 2484 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 0
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_29
timestamp 0
transform 1 0 3772 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_41
timestamp 0
transform 1 0 4876 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_53
timestamp 0
transform 1 0 5980 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_65
timestamp 0
transform 1 0 7084 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_77
timestamp 0
transform 1 0 8188 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_83
timestamp 0
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_85
timestamp 0
transform 1 0 8924 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_97
timestamp 0
transform 1 0 10028 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_109
timestamp 0
transform 1 0 11132 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_121
timestamp 0
transform 1 0 12236 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 0
transform 1 0 13340 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 0
transform 1 0 13892 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 0
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 0
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 0
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_177
timestamp 0
transform 1 0 17388 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_189
timestamp 0
transform 1 0 18492 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 0
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_197
timestamp 0
transform 1 0 19228 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_209
timestamp 0
transform 1 0 20332 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_213
timestamp 0
transform 1 0 20700 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_234
timestamp 0
transform 1 0 22632 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_248
timestamp 0
transform 1 0 23920 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_260
timestamp 0
transform 1 0 25024 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_303
timestamp 0
transform 1 0 28980 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_307
timestamp 0
transform 1 0 29348 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_317
timestamp 0
transform 1 0 30268 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_329
timestamp 0
transform 1 0 31372 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_341
timestamp 0
transform 1 0 32476 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_353
timestamp 0
transform 1 0 33580 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_361
timestamp 0
transform 1 0 34316 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_365
timestamp 0
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_377
timestamp 0
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_389
timestamp 0
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_401
timestamp 0
transform 1 0 37996 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_3
timestamp 0
transform 1 0 1380 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_15
timestamp 0
transform 1 0 2484 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_27
timestamp 0
transform 1 0 3588 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_39
timestamp 0
transform 1 0 4692 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_51
timestamp 0
transform 1 0 5796 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_55
timestamp 0
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_57
timestamp 0
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_69
timestamp 0
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_81
timestamp 0
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_93
timestamp 0
transform 1 0 9660 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_105
timestamp 0
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 0
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 0
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 0
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_137
timestamp 0
transform 1 0 13708 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_149
timestamp 0
transform 1 0 14812 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_161
timestamp 0
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_167
timestamp 0
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_169
timestamp 0
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_181
timestamp 0
transform 1 0 17756 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_193
timestamp 0
transform 1 0 18860 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_205
timestamp 0
transform 1 0 19964 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_217
timestamp 0
transform 1 0 21068 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_222
timestamp 0
transform 1 0 21528 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_253
timestamp 0
transform 1 0 24380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_278
timestamp 0
transform 1 0 26680 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_289
timestamp 0
transform 1 0 27692 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_310
timestamp 0
transform 1 0 29624 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_322
timestamp 0
transform 1 0 30728 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_334
timestamp 0
transform 1 0 31832 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_337
timestamp 0
transform 1 0 32108 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_349
timestamp 0
transform 1 0 33212 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_361
timestamp 0
transform 1 0 34316 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_373
timestamp 0
transform 1 0 35420 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_385
timestamp 0
transform 1 0 36524 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_391
timestamp 0
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_393
timestamp 0
transform 1 0 37260 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_405
timestamp 0
transform 1 0 38364 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_3
timestamp 0
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_15
timestamp 0
transform 1 0 2484 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 0
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_29
timestamp 0
transform 1 0 3772 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_41
timestamp 0
transform 1 0 4876 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_53
timestamp 0
transform 1 0 5980 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_65
timestamp 0
transform 1 0 7084 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_77
timestamp 0
transform 1 0 8188 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_83
timestamp 0
transform 1 0 8740 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_85
timestamp 0
transform 1 0 8924 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_97
timestamp 0
transform 1 0 10028 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_109
timestamp 0
transform 1 0 11132 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_121
timestamp 0
transform 1 0 12236 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_133
timestamp 0
transform 1 0 13340 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_139
timestamp 0
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_141
timestamp 0
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_153
timestamp 0
transform 1 0 15180 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_165
timestamp 0
transform 1 0 16284 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_177
timestamp 0
transform 1 0 17388 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_189
timestamp 0
transform 1 0 18492 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 0
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_197
timestamp 0
transform 1 0 19228 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_209
timestamp 0
transform 1 0 20332 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_262
timestamp 0
transform 1 0 25208 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_305
timestamp 0
transform 1 0 29164 0 1 10880
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_315
timestamp 0
transform 1 0 30084 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_327
timestamp 0
transform 1 0 31188 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_339
timestamp 0
transform 1 0 32292 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_351
timestamp 0
transform 1 0 33396 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_363
timestamp 0
transform 1 0 34500 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_365
timestamp 0
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_377
timestamp 0
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_389
timestamp 0
transform 1 0 36892 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_401
timestamp 0
transform 1 0 37996 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_3
timestamp 0
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_15
timestamp 0
transform 1 0 2484 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_27
timestamp 0
transform 1 0 3588 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_39
timestamp 0
transform 1 0 4692 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_51
timestamp 0
transform 1 0 5796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 0
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 0
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 0
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 0
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_93
timestamp 0
transform 1 0 9660 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_105
timestamp 0
transform 1 0 10764 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_111
timestamp 0
transform 1 0 11316 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 0
transform 1 0 11500 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_125
timestamp 0
transform 1 0 12604 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_137
timestamp 0
transform 1 0 13708 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_149
timestamp 0
transform 1 0 14812 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 0
transform 1 0 15916 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 0
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 0
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_181
timestamp 0
transform 1 0 17756 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_189
timestamp 0
transform 1 0 18492 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_217
timestamp 0
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 0
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_237
timestamp 0
transform 1 0 22908 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_270
timestamp 0
transform 1 0 25944 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_286
timestamp 0
transform 1 0 27416 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_314
timestamp 0
transform 1 0 29992 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_326
timestamp 0
transform 1 0 31096 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_334
timestamp 0
transform 1 0 31832 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_337
timestamp 0
transform 1 0 32108 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_349
timestamp 0
transform 1 0 33212 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_361
timestamp 0
transform 1 0 34316 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_373
timestamp 0
transform 1 0 35420 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_385
timestamp 0
transform 1 0 36524 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_391
timestamp 0
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_393
timestamp 0
transform 1 0 37260 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_405
timestamp 0
transform 1 0 38364 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_3
timestamp 0
transform 1 0 1380 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_15
timestamp 0
transform 1 0 2484 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_27
timestamp 0
transform 1 0 3588 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_29
timestamp 0
transform 1 0 3772 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_41
timestamp 0
transform 1 0 4876 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_53
timestamp 0
transform 1 0 5980 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_65
timestamp 0
transform 1 0 7084 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_77
timestamp 0
transform 1 0 8188 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 0
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_85
timestamp 0
transform 1 0 8924 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_97
timestamp 0
transform 1 0 10028 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_109
timestamp 0
transform 1 0 11132 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_121
timestamp 0
transform 1 0 12236 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_133
timestamp 0
transform 1 0 13340 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_139
timestamp 0
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 0
transform 1 0 14076 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_153
timestamp 0
transform 1 0 15180 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_165
timestamp 0
transform 1 0 16284 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_177
timestamp 0
transform 1 0 17388 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_183
timestamp 0
transform 1 0 17940 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_217
timestamp 0
transform 1 0 21068 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_221
timestamp 0
transform 1 0 21436 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_239
timestamp 0
transform 1 0 23092 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_253
timestamp 0
transform 1 0 24380 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_260
timestamp 0
transform 1 0 25024 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_278
timestamp 0
transform 1 0 26680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_290
timestamp 0
transform 1 0 27784 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_295
timestamp 0
transform 1 0 28244 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_307
timestamp 0
transform 1 0 29348 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_309
timestamp 0
transform 1 0 29532 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_321
timestamp 0
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_333
timestamp 0
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_345
timestamp 0
transform 1 0 32844 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_357
timestamp 0
transform 1 0 33948 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_363
timestamp 0
transform 1 0 34500 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_365
timestamp 0
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_377
timestamp 0
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_389
timestamp 0
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_401
timestamp 0
transform 1 0 37996 0 1 11968
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_6
timestamp 0
transform 1 0 1656 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_18
timestamp 0
transform 1 0 2760 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_30
timestamp 0
transform 1 0 3864 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_42
timestamp 0
transform 1 0 4968 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_54
timestamp 0
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_57
timestamp 0
transform 1 0 6348 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_69
timestamp 0
transform 1 0 7452 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_81
timestamp 0
transform 1 0 8556 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_93
timestamp 0
transform 1 0 9660 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_105
timestamp 0
transform 1 0 10764 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_111
timestamp 0
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_113
timestamp 0
transform 1 0 11500 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_125
timestamp 0
transform 1 0 12604 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_137
timestamp 0
transform 1 0 13708 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_149
timestamp 0
transform 1 0 14812 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_161
timestamp 0
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 0
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_169
timestamp 0
transform 1 0 16652 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_181
timestamp 0
transform 1 0 17756 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_193
timestamp 0
transform 1 0 18860 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_208
timestamp 0
transform 1 0 20240 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_218
timestamp 0
transform 1 0 21160 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_222
timestamp 0
transform 1 0 21528 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_274
timestamp 0
transform 1 0 26312 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_281
timestamp 0
transform 1 0 26956 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_285
timestamp 0
transform 1 0 27324 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_309
timestamp 0
transform 1 0 29532 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_321
timestamp 0
transform 1 0 30636 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_333
timestamp 0
transform 1 0 31740 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_337
timestamp 0
transform 1 0 32108 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_349
timestamp 0
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_361
timestamp 0
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_373
timestamp 0
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_385
timestamp 0
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_391
timestamp 0
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_393
timestamp 0
transform 1 0 37260 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_405
timestamp 0
transform 1 0 38364 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 0
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 0
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 0
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_29
timestamp 0
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_41
timestamp 0
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_53
timestamp 0
transform 1 0 5980 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_65
timestamp 0
transform 1 0 7084 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_77
timestamp 0
transform 1 0 8188 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_83
timestamp 0
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_85
timestamp 0
transform 1 0 8924 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_97
timestamp 0
transform 1 0 10028 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_109
timestamp 0
transform 1 0 11132 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_121
timestamp 0
transform 1 0 12236 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_133
timestamp 0
transform 1 0 13340 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 0
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_141
timestamp 0
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_153
timestamp 0
transform 1 0 15180 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_165
timestamp 0
transform 1 0 16284 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_177
timestamp 0
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_189
timestamp 0
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_195
timestamp 0
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_204
timestamp 0
transform 1 0 19872 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_235
timestamp 0
transform 1 0 22724 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_239
timestamp 0
transform 1 0 23092 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_253
timestamp 0
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_257
timestamp 0
transform 1 0 24748 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_297
timestamp 0
transform 1 0 28428 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_20_305
timestamp 0
transform 1 0 29164 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_309
timestamp 0
transform 1 0 29532 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_321
timestamp 0
transform 1 0 30636 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_333
timestamp 0
transform 1 0 31740 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_345
timestamp 0
transform 1 0 32844 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_357
timestamp 0
transform 1 0 33948 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_363
timestamp 0
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_365
timestamp 0
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_377
timestamp 0
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_389
timestamp 0
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_401
timestamp 0
transform 1 0 37996 0 1 13056
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_3
timestamp 0
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_15
timestamp 0
transform 1 0 2484 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_27
timestamp 0
transform 1 0 3588 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_39
timestamp 0
transform 1 0 4692 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_51
timestamp 0
transform 1 0 5796 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_55
timestamp 0
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_57
timestamp 0
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_69
timestamp 0
transform 1 0 7452 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_81
timestamp 0
transform 1 0 8556 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_93
timestamp 0
transform 1 0 9660 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_105
timestamp 0
transform 1 0 10764 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 0
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 0
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 0
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_137
timestamp 0
transform 1 0 13708 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_149
timestamp 0
transform 1 0 14812 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 0
transform 1 0 15916 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 0
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_169
timestamp 0
transform 1 0 16652 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_181
timestamp 0
transform 1 0 17756 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_189
timestamp 0
transform 1 0 18492 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_218
timestamp 0
transform 1 0 21160 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_232
timestamp 0
transform 1 0 22448 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_236
timestamp 0
transform 1 0 22816 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_257
timestamp 0
transform 1 0 24748 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_278
timestamp 0
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_292
timestamp 0
transform 1 0 27968 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_304
timestamp 0
transform 1 0 29072 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_316
timestamp 0
transform 1 0 30176 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_328
timestamp 0
transform 1 0 31280 0 -1 14144
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_337
timestamp 0
transform 1 0 32108 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_349
timestamp 0
transform 1 0 33212 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_361
timestamp 0
transform 1 0 34316 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_373
timestamp 0
transform 1 0 35420 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_385
timestamp 0
transform 1 0 36524 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_391
timestamp 0
transform 1 0 37076 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_393
timestamp 0
transform 1 0 37260 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_405
timestamp 0
transform 1 0 38364 0 -1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_3
timestamp 0
transform 1 0 1380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_15
timestamp 0
transform 1 0 2484 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 0
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_29
timestamp 0
transform 1 0 3772 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_41
timestamp 0
transform 1 0 4876 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_53
timestamp 0
transform 1 0 5980 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_65
timestamp 0
transform 1 0 7084 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_77
timestamp 0
transform 1 0 8188 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_83
timestamp 0
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_85
timestamp 0
transform 1 0 8924 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_97
timestamp 0
transform 1 0 10028 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_109
timestamp 0
transform 1 0 11132 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_121
timestamp 0
transform 1 0 12236 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_133
timestamp 0
transform 1 0 13340 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 0
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 0
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_153
timestamp 0
transform 1 0 15180 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_165
timestamp 0
transform 1 0 16284 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_177
timestamp 0
transform 1 0 17388 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_189
timestamp 0
transform 1 0 18492 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 0
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_206
timestamp 0
transform 1 0 20056 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_261
timestamp 0
transform 1 0 25116 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_295
timestamp 0
transform 1 0 28244 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 0
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_309
timestamp 0
transform 1 0 29532 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_321
timestamp 0
transform 1 0 30636 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_333
timestamp 0
transform 1 0 31740 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_345
timestamp 0
transform 1 0 32844 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_357
timestamp 0
transform 1 0 33948 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_363
timestamp 0
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_365
timestamp 0
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_377
timestamp 0
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_389
timestamp 0
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_401
timestamp 0
transform 1 0 37996 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 0
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_15
timestamp 0
transform 1 0 2484 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_27
timestamp 0
transform 1 0 3588 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_39
timestamp 0
transform 1 0 4692 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_51
timestamp 0
transform 1 0 5796 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_55
timestamp 0
transform 1 0 6164 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_57
timestamp 0
transform 1 0 6348 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_69
timestamp 0
transform 1 0 7452 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_81
timestamp 0
transform 1 0 8556 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_93
timestamp 0
transform 1 0 9660 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_105
timestamp 0
transform 1 0 10764 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 0
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_113
timestamp 0
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_125
timestamp 0
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_137
timestamp 0
transform 1 0 13708 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_149
timestamp 0
transform 1 0 14812 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_161
timestamp 0
transform 1 0 15916 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_167
timestamp 0
transform 1 0 16468 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_169
timestamp 0
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_181
timestamp 0
transform 1 0 17756 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_189
timestamp 0
transform 1 0 18492 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_195
timestamp 0
transform 1 0 19044 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_203
timestamp 0
transform 1 0 19780 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_234
timestamp 0
transform 1 0 22632 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_240
timestamp 0
transform 1 0 23184 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_268
timestamp 0
transform 1 0 25760 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_281
timestamp 0
transform 1 0 26956 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_293
timestamp 0
transform 1 0 28060 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_305
timestamp 0
transform 1 0 29164 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_317
timestamp 0
transform 1 0 30268 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_329
timestamp 0
transform 1 0 31372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_335
timestamp 0
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_337
timestamp 0
transform 1 0 32108 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_349
timestamp 0
transform 1 0 33212 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_361
timestamp 0
transform 1 0 34316 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_373
timestamp 0
transform 1 0 35420 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_385
timestamp 0
transform 1 0 36524 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_391
timestamp 0
transform 1 0 37076 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_393
timestamp 0
transform 1 0 37260 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_405
timestamp 0
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_3
timestamp 0
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_15
timestamp 0
transform 1 0 2484 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 0
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_29
timestamp 0
transform 1 0 3772 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_41
timestamp 0
transform 1 0 4876 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_53
timestamp 0
transform 1 0 5980 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_65
timestamp 0
transform 1 0 7084 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_77
timestamp 0
transform 1 0 8188 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 0
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_85
timestamp 0
transform 1 0 8924 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_97
timestamp 0
transform 1 0 10028 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_109
timestamp 0
transform 1 0 11132 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_121
timestamp 0
transform 1 0 12236 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_133
timestamp 0
transform 1 0 13340 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_139
timestamp 0
transform 1 0 13892 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_141
timestamp 0
transform 1 0 14076 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_153
timestamp 0
transform 1 0 15180 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_165
timestamp 0
transform 1 0 16284 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_177
timestamp 0
transform 1 0 17388 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_189
timestamp 0
transform 1 0 18492 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 0
transform 1 0 19044 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_197
timestamp 0
transform 1 0 19228 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_209
timestamp 0
transform 1 0 20332 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_214
timestamp 0
transform 1 0 20792 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_221
timestamp 0
transform 1 0 21436 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_247
timestamp 0
transform 1 0 23828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 0
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_260
timestamp 0
transform 1 0 25024 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_272
timestamp 0
transform 1 0 26128 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_284
timestamp 0
transform 1 0 27232 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_296
timestamp 0
transform 1 0 28336 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_309
timestamp 0
transform 1 0 29532 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_321
timestamp 0
transform 1 0 30636 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_333
timestamp 0
transform 1 0 31740 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_345
timestamp 0
transform 1 0 32844 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_357
timestamp 0
transform 1 0 33948 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_363
timestamp 0
transform 1 0 34500 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_365
timestamp 0
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_377
timestamp 0
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_389
timestamp 0
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_401
timestamp 0
transform 1 0 37996 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_3
timestamp 0
transform 1 0 1380 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_15
timestamp 0
transform 1 0 2484 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_27
timestamp 0
transform 1 0 3588 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_39
timestamp 0
transform 1 0 4692 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_51
timestamp 0
transform 1 0 5796 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_55
timestamp 0
transform 1 0 6164 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 0
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 0
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_81
timestamp 0
transform 1 0 8556 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_93
timestamp 0
transform 1 0 9660 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_105
timestamp 0
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 0
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 0
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 0
transform 1 0 12604 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_137
timestamp 0
transform 1 0 13708 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 0
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 0
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 0
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 0
transform 1 0 16652 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_181
timestamp 0
transform 1 0 17756 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_193
timestamp 0
transform 1 0 18860 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_205
timestamp 0
transform 1 0 19964 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_217
timestamp 0
transform 1 0 21068 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 0
transform 1 0 21620 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_225
timestamp 0
transform 1 0 21804 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_229
timestamp 0
transform 1 0 22172 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_238
timestamp 0
transform 1 0 23000 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_242
timestamp 0
transform 1 0 23368 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_250
timestamp 0
transform 1 0 24104 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_262
timestamp 0
transform 1 0 25208 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_274
timestamp 0
transform 1 0 26312 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_281
timestamp 0
transform 1 0 26956 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_293
timestamp 0
transform 1 0 28060 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_305
timestamp 0
transform 1 0 29164 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_317
timestamp 0
transform 1 0 30268 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_329
timestamp 0
transform 1 0 31372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_335
timestamp 0
transform 1 0 31924 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_337
timestamp 0
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_349
timestamp 0
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_361
timestamp 0
transform 1 0 34316 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_373
timestamp 0
transform 1 0 35420 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_385
timestamp 0
transform 1 0 36524 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_391
timestamp 0
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_393
timestamp 0
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_405
timestamp 0
transform 1 0 38364 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_3
timestamp 0
transform 1 0 1380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_15
timestamp 0
transform 1 0 2484 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 0
transform 1 0 3588 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_29
timestamp 0
transform 1 0 3772 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_41
timestamp 0
transform 1 0 4876 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_53
timestamp 0
transform 1 0 5980 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_65
timestamp 0
transform 1 0 7084 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_77
timestamp 0
transform 1 0 8188 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_83
timestamp 0
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_85
timestamp 0
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_97
timestamp 0
transform 1 0 10028 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_109
timestamp 0
transform 1 0 11132 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_121
timestamp 0
transform 1 0 12236 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_133
timestamp 0
transform 1 0 13340 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 0
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_141
timestamp 0
transform 1 0 14076 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_153
timestamp 0
transform 1 0 15180 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_165
timestamp 0
transform 1 0 16284 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_177
timestamp 0
transform 1 0 17388 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_189
timestamp 0
transform 1 0 18492 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_195
timestamp 0
transform 1 0 19044 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_197
timestamp 0
transform 1 0 19228 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_209
timestamp 0
transform 1 0 20332 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_221
timestamp 0
transform 1 0 21436 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_233
timestamp 0
transform 1 0 22540 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_245
timestamp 0
transform 1 0 23644 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_251
timestamp 0
transform 1 0 24196 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_253
timestamp 0
transform 1 0 24380 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_265
timestamp 0
transform 1 0 25484 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_277
timestamp 0
transform 1 0 26588 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_289
timestamp 0
transform 1 0 27692 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_301
timestamp 0
transform 1 0 28796 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_307
timestamp 0
transform 1 0 29348 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_309
timestamp 0
transform 1 0 29532 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_321
timestamp 0
transform 1 0 30636 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_333
timestamp 0
transform 1 0 31740 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_345
timestamp 0
transform 1 0 32844 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_357
timestamp 0
transform 1 0 33948 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_363
timestamp 0
transform 1 0 34500 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_365
timestamp 0
transform 1 0 34684 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_377
timestamp 0
transform 1 0 35788 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_389
timestamp 0
transform 1 0 36892 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_401
timestamp 0
transform 1 0 37996 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 0
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_15
timestamp 0
transform 1 0 2484 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_27
timestamp 0
transform 1 0 3588 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_39
timestamp 0
transform 1 0 4692 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_51
timestamp 0
transform 1 0 5796 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 0
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 0
transform 1 0 6348 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_69
timestamp 0
transform 1 0 7452 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_81
timestamp 0
transform 1 0 8556 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_93
timestamp 0
transform 1 0 9660 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_105
timestamp 0
transform 1 0 10764 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_111
timestamp 0
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_113
timestamp 0
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_125
timestamp 0
transform 1 0 12604 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_137
timestamp 0
transform 1 0 13708 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_149
timestamp 0
transform 1 0 14812 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_161
timestamp 0
transform 1 0 15916 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 0
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_169
timestamp 0
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_181
timestamp 0
transform 1 0 17756 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_193
timestamp 0
transform 1 0 18860 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_205
timestamp 0
transform 1 0 19964 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_217
timestamp 0
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 0
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_225
timestamp 0
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_237
timestamp 0
transform 1 0 22908 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_249
timestamp 0
transform 1 0 24012 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_261
timestamp 0
transform 1 0 25116 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_273
timestamp 0
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_279
timestamp 0
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_281
timestamp 0
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_293
timestamp 0
transform 1 0 28060 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_305
timestamp 0
transform 1 0 29164 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_317
timestamp 0
transform 1 0 30268 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_329
timestamp 0
transform 1 0 31372 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_335
timestamp 0
transform 1 0 31924 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_337
timestamp 0
transform 1 0 32108 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_349
timestamp 0
transform 1 0 33212 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_361
timestamp 0
transform 1 0 34316 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_373
timestamp 0
transform 1 0 35420 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_385
timestamp 0
transform 1 0 36524 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_391
timestamp 0
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_393
timestamp 0
transform 1 0 37260 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_405
timestamp 0
transform 1 0 38364 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_3
timestamp 0
transform 1 0 1380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_15
timestamp 0
transform 1 0 2484 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_27
timestamp 0
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_29
timestamp 0
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_41
timestamp 0
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_53
timestamp 0
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_65
timestamp 0
transform 1 0 7084 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_77
timestamp 0
transform 1 0 8188 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_83
timestamp 0
transform 1 0 8740 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 0
transform 1 0 8924 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_97
timestamp 0
transform 1 0 10028 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_109
timestamp 0
transform 1 0 11132 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_121
timestamp 0
transform 1 0 12236 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_133
timestamp 0
transform 1 0 13340 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_139
timestamp 0
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_141
timestamp 0
transform 1 0 14076 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_153
timestamp 0
transform 1 0 15180 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_165
timestamp 0
transform 1 0 16284 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_177
timestamp 0
transform 1 0 17388 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_189
timestamp 0
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 0
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 0
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_209
timestamp 0
transform 1 0 20332 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_221
timestamp 0
transform 1 0 21436 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_233
timestamp 0
transform 1 0 22540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_245
timestamp 0
transform 1 0 23644 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_251
timestamp 0
transform 1 0 24196 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_253
timestamp 0
transform 1 0 24380 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_265
timestamp 0
transform 1 0 25484 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_277
timestamp 0
transform 1 0 26588 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_289
timestamp 0
transform 1 0 27692 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_301
timestamp 0
transform 1 0 28796 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_307
timestamp 0
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_309
timestamp 0
transform 1 0 29532 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_321
timestamp 0
transform 1 0 30636 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_333
timestamp 0
transform 1 0 31740 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_345
timestamp 0
transform 1 0 32844 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_357
timestamp 0
transform 1 0 33948 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_363
timestamp 0
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_365
timestamp 0
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_377
timestamp 0
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_389
timestamp 0
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_401
timestamp 0
transform 1 0 37996 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_3
timestamp 0
transform 1 0 1380 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_15
timestamp 0
transform 1 0 2484 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_27
timestamp 0
transform 1 0 3588 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_39
timestamp 0
transform 1 0 4692 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_51
timestamp 0
transform 1 0 5796 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_55
timestamp 0
transform 1 0 6164 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 0
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_69
timestamp 0
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_81
timestamp 0
transform 1 0 8556 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_93
timestamp 0
transform 1 0 9660 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_105
timestamp 0
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 0
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_113
timestamp 0
transform 1 0 11500 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 0
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_137
timestamp 0
transform 1 0 13708 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_149
timestamp 0
transform 1 0 14812 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_161
timestamp 0
transform 1 0 15916 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 0
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_169
timestamp 0
transform 1 0 16652 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_181
timestamp 0
transform 1 0 17756 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_193
timestamp 0
transform 1 0 18860 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_205
timestamp 0
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_217
timestamp 0
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 0
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_225
timestamp 0
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_237
timestamp 0
transform 1 0 22908 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_249
timestamp 0
transform 1 0 24012 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_261
timestamp 0
transform 1 0 25116 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_273
timestamp 0
transform 1 0 26220 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_279
timestamp 0
transform 1 0 26772 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_281
timestamp 0
transform 1 0 26956 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_293
timestamp 0
transform 1 0 28060 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_305
timestamp 0
transform 1 0 29164 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_317
timestamp 0
transform 1 0 30268 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_329
timestamp 0
transform 1 0 31372 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_335
timestamp 0
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_337
timestamp 0
transform 1 0 32108 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_349
timestamp 0
transform 1 0 33212 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_361
timestamp 0
transform 1 0 34316 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_373
timestamp 0
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_385
timestamp 0
transform 1 0 36524 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_391
timestamp 0
transform 1 0 37076 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_393
timestamp 0
transform 1 0 37260 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_405
timestamp 0
transform 1 0 38364 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_3
timestamp 0
transform 1 0 1380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_15
timestamp 0
transform 1 0 2484 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_27
timestamp 0
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_29
timestamp 0
transform 1 0 3772 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 0
transform 1 0 4876 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 0
transform 1 0 5980 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_65
timestamp 0
transform 1 0 7084 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_77
timestamp 0
transform 1 0 8188 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_83
timestamp 0
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 0
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_97
timestamp 0
transform 1 0 10028 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_109
timestamp 0
transform 1 0 11132 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 0
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 0
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 0
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_141
timestamp 0
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_153
timestamp 0
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_165
timestamp 0
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_177
timestamp 0
transform 1 0 17388 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_189
timestamp 0
transform 1 0 18492 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 0
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_197
timestamp 0
transform 1 0 19228 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_209
timestamp 0
transform 1 0 20332 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_221
timestamp 0
transform 1 0 21436 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_233
timestamp 0
transform 1 0 22540 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_245
timestamp 0
transform 1 0 23644 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 0
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 0
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 0
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 0
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_289
timestamp 0
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_301
timestamp 0
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 0
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 0
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_321
timestamp 0
transform 1 0 30636 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_333
timestamp 0
transform 1 0 31740 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_345
timestamp 0
transform 1 0 32844 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_357
timestamp 0
transform 1 0 33948 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_363
timestamp 0
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_365
timestamp 0
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_377
timestamp 0
transform 1 0 35788 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_389
timestamp 0
transform 1 0 36892 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_401
timestamp 0
transform 1 0 37996 0 1 18496
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_3
timestamp 0
transform 1 0 1380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_15
timestamp 0
transform 1 0 2484 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_27
timestamp 0
transform 1 0 3588 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_39
timestamp 0
transform 1 0 4692 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_51
timestamp 0
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_55
timestamp 0
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 0
transform 1 0 6348 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 0
transform 1 0 7452 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_81
timestamp 0
transform 1 0 8556 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_93
timestamp 0
transform 1 0 9660 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 0
transform 1 0 10764 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 0
transform 1 0 11316 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_113
timestamp 0
transform 1 0 11500 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_125
timestamp 0
transform 1 0 12604 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_137
timestamp 0
transform 1 0 13708 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_149
timestamp 0
transform 1 0 14812 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_161
timestamp 0
transform 1 0 15916 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_167
timestamp 0
transform 1 0 16468 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_169
timestamp 0
transform 1 0 16652 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_181
timestamp 0
transform 1 0 17756 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_193
timestamp 0
transform 1 0 18860 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_205
timestamp 0
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 0
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 0
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_225
timestamp 0
transform 1 0 21804 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_237
timestamp 0
transform 1 0 22908 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_249
timestamp 0
transform 1 0 24012 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_261
timestamp 0
transform 1 0 25116 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_273
timestamp 0
transform 1 0 26220 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_279
timestamp 0
transform 1 0 26772 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_281
timestamp 0
transform 1 0 26956 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_293
timestamp 0
transform 1 0 28060 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_305
timestamp 0
transform 1 0 29164 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_317
timestamp 0
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_329
timestamp 0
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_335
timestamp 0
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_337
timestamp 0
transform 1 0 32108 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_349
timestamp 0
transform 1 0 33212 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_361
timestamp 0
transform 1 0 34316 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_373
timestamp 0
transform 1 0 35420 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_385
timestamp 0
transform 1 0 36524 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_391
timestamp 0
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_393
timestamp 0
transform 1 0 37260 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_405
timestamp 0
transform 1 0 38364 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_3
timestamp 0
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_15
timestamp 0
transform 1 0 2484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 0
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_29
timestamp 0
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_41
timestamp 0
transform 1 0 4876 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_53
timestamp 0
transform 1 0 5980 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_65
timestamp 0
transform 1 0 7084 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_77
timestamp 0
transform 1 0 8188 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 0
transform 1 0 8740 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_85
timestamp 0
transform 1 0 8924 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_97
timestamp 0
transform 1 0 10028 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_109
timestamp 0
transform 1 0 11132 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 0
transform 1 0 12236 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 0
transform 1 0 13340 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 0
transform 1 0 13892 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 0
transform 1 0 14076 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 0
transform 1 0 15180 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_165
timestamp 0
transform 1 0 16284 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_177
timestamp 0
transform 1 0 17388 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_189
timestamp 0
transform 1 0 18492 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 0
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_197
timestamp 0
transform 1 0 19228 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_209
timestamp 0
transform 1 0 20332 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_221
timestamp 0
transform 1 0 21436 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_233
timestamp 0
transform 1 0 22540 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_245
timestamp 0
transform 1 0 23644 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 0
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_253
timestamp 0
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_265
timestamp 0
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_277
timestamp 0
transform 1 0 26588 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_289
timestamp 0
transform 1 0 27692 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_301
timestamp 0
transform 1 0 28796 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_307
timestamp 0
transform 1 0 29348 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_309
timestamp 0
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_321
timestamp 0
transform 1 0 30636 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_333
timestamp 0
transform 1 0 31740 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_345
timestamp 0
transform 1 0 32844 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_357
timestamp 0
transform 1 0 33948 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_363
timestamp 0
transform 1 0 34500 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_365
timestamp 0
transform 1 0 34684 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_377
timestamp 0
transform 1 0 35788 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_389
timestamp 0
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_401
timestamp 0
transform 1 0 37996 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_3
timestamp 0
transform 1 0 1380 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_15
timestamp 0
transform 1 0 2484 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_27
timestamp 0
transform 1 0 3588 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_39
timestamp 0
transform 1 0 4692 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_51
timestamp 0
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_55
timestamp 0
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_57
timestamp 0
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_69
timestamp 0
transform 1 0 7452 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_81
timestamp 0
transform 1 0 8556 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_93
timestamp 0
transform 1 0 9660 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_105
timestamp 0
transform 1 0 10764 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 0
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_113
timestamp 0
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_125
timestamp 0
transform 1 0 12604 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_137
timestamp 0
transform 1 0 13708 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_149
timestamp 0
transform 1 0 14812 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_161
timestamp 0
transform 1 0 15916 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_167
timestamp 0
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_169
timestamp 0
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_181
timestamp 0
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_193
timestamp 0
transform 1 0 18860 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_205
timestamp 0
transform 1 0 19964 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_217
timestamp 0
transform 1 0 21068 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_223
timestamp 0
transform 1 0 21620 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 0
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_237
timestamp 0
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_249
timestamp 0
transform 1 0 24012 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_261
timestamp 0
transform 1 0 25116 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_273
timestamp 0
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_279
timestamp 0
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_281
timestamp 0
transform 1 0 26956 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_293
timestamp 0
transform 1 0 28060 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_305
timestamp 0
transform 1 0 29164 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_317
timestamp 0
transform 1 0 30268 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_329
timestamp 0
transform 1 0 31372 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_335
timestamp 0
transform 1 0 31924 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_337
timestamp 0
transform 1 0 32108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_349
timestamp 0
transform 1 0 33212 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_361
timestamp 0
transform 1 0 34316 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_373
timestamp 0
transform 1 0 35420 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_385
timestamp 0
transform 1 0 36524 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_391
timestamp 0
transform 1 0 37076 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_393
timestamp 0
transform 1 0 37260 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_405
timestamp 0
transform 1 0 38364 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_3
timestamp 0
transform 1 0 1380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_15
timestamp 0
transform 1 0 2484 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 0
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 0
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_41
timestamp 0
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_53
timestamp 0
transform 1 0 5980 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_65
timestamp 0
transform 1 0 7084 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_77
timestamp 0
transform 1 0 8188 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 0
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_85
timestamp 0
transform 1 0 8924 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_97
timestamp 0
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_109
timestamp 0
transform 1 0 11132 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_121
timestamp 0
transform 1 0 12236 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_133
timestamp 0
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 0
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_141
timestamp 0
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_153
timestamp 0
transform 1 0 15180 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_165
timestamp 0
transform 1 0 16284 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_177
timestamp 0
transform 1 0 17388 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_189
timestamp 0
transform 1 0 18492 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_195
timestamp 0
transform 1 0 19044 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_197
timestamp 0
transform 1 0 19228 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_209
timestamp 0
transform 1 0 20332 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_221
timestamp 0
transform 1 0 21436 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_233
timestamp 0
transform 1 0 22540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_245
timestamp 0
transform 1 0 23644 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_251
timestamp 0
transform 1 0 24196 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_253
timestamp 0
transform 1 0 24380 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_265
timestamp 0
transform 1 0 25484 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_277
timestamp 0
transform 1 0 26588 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_289
timestamp 0
transform 1 0 27692 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_301
timestamp 0
transform 1 0 28796 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_307
timestamp 0
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_309
timestamp 0
transform 1 0 29532 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_321
timestamp 0
transform 1 0 30636 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_333
timestamp 0
transform 1 0 31740 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_345
timestamp 0
transform 1 0 32844 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_357
timestamp 0
transform 1 0 33948 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_363
timestamp 0
transform 1 0 34500 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_365
timestamp 0
transform 1 0 34684 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_377
timestamp 0
transform 1 0 35788 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_389
timestamp 0
transform 1 0 36892 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_401
timestamp 0
transform 1 0 37996 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_3
timestamp 0
transform 1 0 1380 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_15
timestamp 0
transform 1 0 2484 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_27
timestamp 0
transform 1 0 3588 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_39
timestamp 0
transform 1 0 4692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 0
transform 1 0 5796 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 0
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 0
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_69
timestamp 0
transform 1 0 7452 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_81
timestamp 0
transform 1 0 8556 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_93
timestamp 0
transform 1 0 9660 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_105
timestamp 0
transform 1 0 10764 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_111
timestamp 0
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_113
timestamp 0
transform 1 0 11500 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_125
timestamp 0
transform 1 0 12604 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_137
timestamp 0
transform 1 0 13708 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_149
timestamp 0
transform 1 0 14812 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_161
timestamp 0
transform 1 0 15916 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 0
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 0
transform 1 0 16652 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_181
timestamp 0
transform 1 0 17756 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_193
timestamp 0
transform 1 0 18860 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_205
timestamp 0
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_217
timestamp 0
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_223
timestamp 0
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_225
timestamp 0
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_237
timestamp 0
transform 1 0 22908 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_249
timestamp 0
transform 1 0 24012 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_261
timestamp 0
transform 1 0 25116 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_273
timestamp 0
transform 1 0 26220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_279
timestamp 0
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_281
timestamp 0
transform 1 0 26956 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_293
timestamp 0
transform 1 0 28060 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_305
timestamp 0
transform 1 0 29164 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_317
timestamp 0
transform 1 0 30268 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_329
timestamp 0
transform 1 0 31372 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_335
timestamp 0
transform 1 0 31924 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_337
timestamp 0
transform 1 0 32108 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_349
timestamp 0
transform 1 0 33212 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_361
timestamp 0
transform 1 0 34316 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_373
timestamp 0
transform 1 0 35420 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_385
timestamp 0
transform 1 0 36524 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_391
timestamp 0
transform 1 0 37076 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_393
timestamp 0
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_405
timestamp 0
transform 1 0 38364 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_3
timestamp 0
transform 1 0 1380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_15
timestamp 0
transform 1 0 2484 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_27
timestamp 0
transform 1 0 3588 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 0
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_41
timestamp 0
transform 1 0 4876 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_53
timestamp 0
transform 1 0 5980 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_65
timestamp 0
transform 1 0 7084 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_77
timestamp 0
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 0
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_85
timestamp 0
transform 1 0 8924 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_97
timestamp 0
transform 1 0 10028 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_109
timestamp 0
transform 1 0 11132 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_121
timestamp 0
transform 1 0 12236 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_133
timestamp 0
transform 1 0 13340 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 0
transform 1 0 13892 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_141
timestamp 0
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_153
timestamp 0
transform 1 0 15180 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_165
timestamp 0
transform 1 0 16284 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_177
timestamp 0
transform 1 0 17388 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_189
timestamp 0
transform 1 0 18492 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_195
timestamp 0
transform 1 0 19044 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_197
timestamp 0
transform 1 0 19228 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_209
timestamp 0
transform 1 0 20332 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_221
timestamp 0
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_233
timestamp 0
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_245
timestamp 0
transform 1 0 23644 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_251
timestamp 0
transform 1 0 24196 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_253
timestamp 0
transform 1 0 24380 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_265
timestamp 0
transform 1 0 25484 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_277
timestamp 0
transform 1 0 26588 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_289
timestamp 0
transform 1 0 27692 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_301
timestamp 0
transform 1 0 28796 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_307
timestamp 0
transform 1 0 29348 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_309
timestamp 0
transform 1 0 29532 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_321
timestamp 0
transform 1 0 30636 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_333
timestamp 0
transform 1 0 31740 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_345
timestamp 0
transform 1 0 32844 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_357
timestamp 0
transform 1 0 33948 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_363
timestamp 0
transform 1 0 34500 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_365
timestamp 0
transform 1 0 34684 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_377
timestamp 0
transform 1 0 35788 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_389
timestamp 0
transform 1 0 36892 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_401
timestamp 0
transform 1 0 37996 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 0
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_15
timestamp 0
transform 1 0 2484 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_27
timestamp 0
transform 1 0 3588 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_39
timestamp 0
transform 1 0 4692 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 0
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 0
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 0
transform 1 0 6348 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_69
timestamp 0
transform 1 0 7452 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_81
timestamp 0
transform 1 0 8556 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_93
timestamp 0
transform 1 0 9660 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_105
timestamp 0
transform 1 0 10764 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 0
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_113
timestamp 0
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_125
timestamp 0
transform 1 0 12604 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_137
timestamp 0
transform 1 0 13708 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_149
timestamp 0
transform 1 0 14812 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_161
timestamp 0
transform 1 0 15916 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 0
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_169
timestamp 0
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_181
timestamp 0
transform 1 0 17756 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_193
timestamp 0
transform 1 0 18860 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_205
timestamp 0
transform 1 0 19964 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_217
timestamp 0
transform 1 0 21068 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 0
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_225
timestamp 0
transform 1 0 21804 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_237
timestamp 0
transform 1 0 22908 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_249
timestamp 0
transform 1 0 24012 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_261
timestamp 0
transform 1 0 25116 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_273
timestamp 0
transform 1 0 26220 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_279
timestamp 0
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_281
timestamp 0
transform 1 0 26956 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_293
timestamp 0
transform 1 0 28060 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_305
timestamp 0
transform 1 0 29164 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_317
timestamp 0
transform 1 0 30268 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_329
timestamp 0
transform 1 0 31372 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_335
timestamp 0
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_337
timestamp 0
transform 1 0 32108 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_349
timestamp 0
transform 1 0 33212 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_361
timestamp 0
transform 1 0 34316 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_373
timestamp 0
transform 1 0 35420 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_385
timestamp 0
transform 1 0 36524 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_391
timestamp 0
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_393
timestamp 0
transform 1 0 37260 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_405
timestamp 0
transform 1 0 38364 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_3
timestamp 0
transform 1 0 1380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_15
timestamp 0
transform 1 0 2484 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_27
timestamp 0
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 0
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_41
timestamp 0
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_53
timestamp 0
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_65
timestamp 0
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 0
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 0
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_85
timestamp 0
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_97
timestamp 0
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_109
timestamp 0
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_121
timestamp 0
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_133
timestamp 0
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_139
timestamp 0
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_141
timestamp 0
transform 1 0 14076 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_153
timestamp 0
transform 1 0 15180 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_165
timestamp 0
transform 1 0 16284 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_177
timestamp 0
transform 1 0 17388 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_189
timestamp 0
transform 1 0 18492 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_195
timestamp 0
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 0
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_209
timestamp 0
transform 1 0 20332 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_221
timestamp 0
transform 1 0 21436 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_233
timestamp 0
transform 1 0 22540 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_245
timestamp 0
transform 1 0 23644 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_251
timestamp 0
transform 1 0 24196 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_253
timestamp 0
transform 1 0 24380 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_265
timestamp 0
transform 1 0 25484 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_277
timestamp 0
transform 1 0 26588 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_289
timestamp 0
transform 1 0 27692 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_301
timestamp 0
transform 1 0 28796 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_307
timestamp 0
transform 1 0 29348 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_309
timestamp 0
transform 1 0 29532 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_321
timestamp 0
transform 1 0 30636 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_333
timestamp 0
transform 1 0 31740 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_345
timestamp 0
transform 1 0 32844 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_357
timestamp 0
transform 1 0 33948 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_363
timestamp 0
transform 1 0 34500 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_365
timestamp 0
transform 1 0 34684 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_377
timestamp 0
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_389
timestamp 0
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_401
timestamp 0
transform 1 0 37996 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 0
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 0
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 0
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_39
timestamp 0
transform 1 0 4692 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_51
timestamp 0
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_55
timestamp 0
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_57
timestamp 0
transform 1 0 6348 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_69
timestamp 0
transform 1 0 7452 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_81
timestamp 0
transform 1 0 8556 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_93
timestamp 0
transform 1 0 9660 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_105
timestamp 0
transform 1 0 10764 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 0
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 0
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_125
timestamp 0
transform 1 0 12604 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_137
timestamp 0
transform 1 0 13708 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_149
timestamp 0
transform 1 0 14812 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_161
timestamp 0
transform 1 0 15916 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 0
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 0
transform 1 0 16652 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_181
timestamp 0
transform 1 0 17756 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_193
timestamp 0
transform 1 0 18860 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_205
timestamp 0
transform 1 0 19964 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_217
timestamp 0
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_223
timestamp 0
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_225
timestamp 0
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_237
timestamp 0
transform 1 0 22908 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_249
timestamp 0
transform 1 0 24012 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_261
timestamp 0
transform 1 0 25116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_273
timestamp 0
transform 1 0 26220 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_279
timestamp 0
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_281
timestamp 0
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_293
timestamp 0
transform 1 0 28060 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_305
timestamp 0
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_317
timestamp 0
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_329
timestamp 0
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_335
timestamp 0
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_337
timestamp 0
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_349
timestamp 0
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_361
timestamp 0
transform 1 0 34316 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_373
timestamp 0
transform 1 0 35420 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_385
timestamp 0
transform 1 0 36524 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_391
timestamp 0
transform 1 0 37076 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_393
timestamp 0
transform 1 0 37260 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_405
timestamp 0
transform 1 0 38364 0 -1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_3
timestamp 0
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_15
timestamp 0
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 0
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 0
transform 1 0 3772 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 0
transform 1 0 4876 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 0
transform 1 0 5980 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_65
timestamp 0
transform 1 0 7084 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 0
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 0
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 0
transform 1 0 8924 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_97
timestamp 0
transform 1 0 10028 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_109
timestamp 0
transform 1 0 11132 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_121
timestamp 0
transform 1 0 12236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_133
timestamp 0
transform 1 0 13340 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 0
transform 1 0 13892 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_141
timestamp 0
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_153
timestamp 0
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_165
timestamp 0
transform 1 0 16284 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_177
timestamp 0
transform 1 0 17388 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_189
timestamp 0
transform 1 0 18492 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_195
timestamp 0
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 0
transform 1 0 19228 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_209
timestamp 0
transform 1 0 20332 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_221
timestamp 0
transform 1 0 21436 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_233
timestamp 0
transform 1 0 22540 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_245
timestamp 0
transform 1 0 23644 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_251
timestamp 0
transform 1 0 24196 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_253
timestamp 0
transform 1 0 24380 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_265
timestamp 0
transform 1 0 25484 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_277
timestamp 0
transform 1 0 26588 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_289
timestamp 0
transform 1 0 27692 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_301
timestamp 0
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_307
timestamp 0
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_309
timestamp 0
transform 1 0 29532 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_321
timestamp 0
transform 1 0 30636 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_333
timestamp 0
transform 1 0 31740 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_345
timestamp 0
transform 1 0 32844 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_357
timestamp 0
transform 1 0 33948 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_363
timestamp 0
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_365
timestamp 0
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_377
timestamp 0
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_389
timestamp 0
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_401
timestamp 0
transform 1 0 37996 0 1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_3
timestamp 0
transform 1 0 1380 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_15
timestamp 0
transform 1 0 2484 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_27
timestamp 0
transform 1 0 3588 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_39
timestamp 0
transform 1 0 4692 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 0
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 0
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_57
timestamp 0
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_69
timestamp 0
transform 1 0 7452 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_81
timestamp 0
transform 1 0 8556 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_93
timestamp 0
transform 1 0 9660 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_105
timestamp 0
transform 1 0 10764 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_111
timestamp 0
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_113
timestamp 0
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_125
timestamp 0
transform 1 0 12604 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_137
timestamp 0
transform 1 0 13708 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_149
timestamp 0
transform 1 0 14812 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_161
timestamp 0
transform 1 0 15916 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_167
timestamp 0
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_169
timestamp 0
transform 1 0 16652 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_181
timestamp 0
transform 1 0 17756 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_193
timestamp 0
transform 1 0 18860 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_205
timestamp 0
transform 1 0 19964 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_217
timestamp 0
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 0
transform 1 0 21620 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 0
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_237
timestamp 0
transform 1 0 22908 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_249
timestamp 0
transform 1 0 24012 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_261
timestamp 0
transform 1 0 25116 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_273
timestamp 0
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 0
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_281
timestamp 0
transform 1 0 26956 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_293
timestamp 0
transform 1 0 28060 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_305
timestamp 0
transform 1 0 29164 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_317
timestamp 0
transform 1 0 30268 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_329
timestamp 0
transform 1 0 31372 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_335
timestamp 0
transform 1 0 31924 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_337
timestamp 0
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_349
timestamp 0
transform 1 0 33212 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_361
timestamp 0
transform 1 0 34316 0 -1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_373
timestamp 0
transform 1 0 35420 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_385
timestamp 0
transform 1 0 36524 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_391
timestamp 0
transform 1 0 37076 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_393
timestamp 0
transform 1 0 37260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_405
timestamp 0
transform 1 0 38364 0 -1 25024
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_7
timestamp 0
transform 1 0 1748 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_19
timestamp 0
transform 1 0 2852 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 0
transform 1 0 3588 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_29
timestamp 0
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_41
timestamp 0
transform 1 0 4876 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_53
timestamp 0
transform 1 0 5980 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_65
timestamp 0
transform 1 0 7084 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_77
timestamp 0
transform 1 0 8188 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 0
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_85
timestamp 0
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_97
timestamp 0
transform 1 0 10028 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_109
timestamp 0
transform 1 0 11132 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_121
timestamp 0
transform 1 0 12236 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_133
timestamp 0
transform 1 0 13340 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 0
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_141
timestamp 0
transform 1 0 14076 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_153
timestamp 0
transform 1 0 15180 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_165
timestamp 0
transform 1 0 16284 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_177
timestamp 0
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_189
timestamp 0
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_195
timestamp 0
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_197
timestamp 0
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_209
timestamp 0
transform 1 0 20332 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_221
timestamp 0
transform 1 0 21436 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_233
timestamp 0
transform 1 0 22540 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_245
timestamp 0
transform 1 0 23644 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_251
timestamp 0
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_253
timestamp 0
transform 1 0 24380 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_265
timestamp 0
transform 1 0 25484 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_277
timestamp 0
transform 1 0 26588 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_289
timestamp 0
transform 1 0 27692 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_301
timestamp 0
transform 1 0 28796 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_307
timestamp 0
transform 1 0 29348 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_309
timestamp 0
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_321
timestamp 0
transform 1 0 30636 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_333
timestamp 0
transform 1 0 31740 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_345
timestamp 0
transform 1 0 32844 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_357
timestamp 0
transform 1 0 33948 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_363
timestamp 0
transform 1 0 34500 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_365
timestamp 0
transform 1 0 34684 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_377
timestamp 0
transform 1 0 35788 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_389
timestamp 0
transform 1 0 36892 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_401
timestamp 0
transform 1 0 37996 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_3
timestamp 0
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_15
timestamp 0
transform 1 0 2484 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_27
timestamp 0
transform 1 0 3588 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_39
timestamp 0
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 0
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 0
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 0
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 0
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_81
timestamp 0
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_93
timestamp 0
transform 1 0 9660 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_105
timestamp 0
transform 1 0 10764 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 0
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 0
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 0
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_137
timestamp 0
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_149
timestamp 0
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_161
timestamp 0
transform 1 0 15916 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 0
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 0
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_181
timestamp 0
transform 1 0 17756 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_193
timestamp 0
transform 1 0 18860 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_205
timestamp 0
transform 1 0 19964 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_217
timestamp 0
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_223
timestamp 0
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_225
timestamp 0
transform 1 0 21804 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_237
timestamp 0
transform 1 0 22908 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_249
timestamp 0
transform 1 0 24012 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_261
timestamp 0
transform 1 0 25116 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_273
timestamp 0
transform 1 0 26220 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_279
timestamp 0
transform 1 0 26772 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 0
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_293
timestamp 0
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_305
timestamp 0
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_317
timestamp 0
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_329
timestamp 0
transform 1 0 31372 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_335
timestamp 0
transform 1 0 31924 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_337
timestamp 0
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_349
timestamp 0
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_361
timestamp 0
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_373
timestamp 0
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_385
timestamp 0
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_391
timestamp 0
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_393
timestamp 0
transform 1 0 37260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_405
timestamp 0
transform 1 0 38364 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 0
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 0
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 0
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 0
transform 1 0 3772 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_41
timestamp 0
transform 1 0 4876 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_53
timestamp 0
transform 1 0 5980 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_65
timestamp 0
transform 1 0 7084 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_77
timestamp 0
transform 1 0 8188 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_83
timestamp 0
transform 1 0 8740 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 0
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_97
timestamp 0
transform 1 0 10028 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_109
timestamp 0
transform 1 0 11132 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_121
timestamp 0
transform 1 0 12236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_133
timestamp 0
transform 1 0 13340 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_139
timestamp 0
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_141
timestamp 0
transform 1 0 14076 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_153
timestamp 0
transform 1 0 15180 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_165
timestamp 0
transform 1 0 16284 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_177
timestamp 0
transform 1 0 17388 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_189
timestamp 0
transform 1 0 18492 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 0
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_197
timestamp 0
transform 1 0 19228 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_209
timestamp 0
transform 1 0 20332 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_221
timestamp 0
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_233
timestamp 0
transform 1 0 22540 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_245
timestamp 0
transform 1 0 23644 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_251
timestamp 0
transform 1 0 24196 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_253
timestamp 0
transform 1 0 24380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_265
timestamp 0
transform 1 0 25484 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_277
timestamp 0
transform 1 0 26588 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_289
timestamp 0
transform 1 0 27692 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_301
timestamp 0
transform 1 0 28796 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_307
timestamp 0
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_309
timestamp 0
transform 1 0 29532 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_321
timestamp 0
transform 1 0 30636 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_333
timestamp 0
transform 1 0 31740 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_345
timestamp 0
transform 1 0 32844 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_357
timestamp 0
transform 1 0 33948 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_363
timestamp 0
transform 1 0 34500 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_365
timestamp 0
transform 1 0 34684 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_377
timestamp 0
transform 1 0 35788 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_389
timestamp 0
transform 1 0 36892 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_401
timestamp 0
transform 1 0 37996 0 1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 0
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 0
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 0
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 0
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 0
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 0
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 0
transform 1 0 6348 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 0
transform 1 0 7452 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 0
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_93
timestamp 0
transform 1 0 9660 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_105
timestamp 0
transform 1 0 10764 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 0
transform 1 0 11316 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_113
timestamp 0
transform 1 0 11500 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_125
timestamp 0
transform 1 0 12604 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_137
timestamp 0
transform 1 0 13708 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_149
timestamp 0
transform 1 0 14812 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_161
timestamp 0
transform 1 0 15916 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 0
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 0
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_181
timestamp 0
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_193
timestamp 0
transform 1 0 18860 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_205
timestamp 0
transform 1 0 19964 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_217
timestamp 0
transform 1 0 21068 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_223
timestamp 0
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_225
timestamp 0
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_237
timestamp 0
transform 1 0 22908 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_249
timestamp 0
transform 1 0 24012 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_261
timestamp 0
transform 1 0 25116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_273
timestamp 0
transform 1 0 26220 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_279
timestamp 0
transform 1 0 26772 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_281
timestamp 0
transform 1 0 26956 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_293
timestamp 0
transform 1 0 28060 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_305
timestamp 0
transform 1 0 29164 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_317
timestamp 0
transform 1 0 30268 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_329
timestamp 0
transform 1 0 31372 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_335
timestamp 0
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_337
timestamp 0
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_349
timestamp 0
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_361
timestamp 0
transform 1 0 34316 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_373
timestamp 0
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_385
timestamp 0
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_391
timestamp 0
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_393
timestamp 0
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_405
timestamp 0
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 0
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 0
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 0
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_29
timestamp 0
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 0
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_53
timestamp 0
transform 1 0 5980 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_65
timestamp 0
transform 1 0 7084 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_77
timestamp 0
transform 1 0 8188 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_83
timestamp 0
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_85
timestamp 0
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_97
timestamp 0
transform 1 0 10028 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_109
timestamp 0
transform 1 0 11132 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_121
timestamp 0
transform 1 0 12236 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_133
timestamp 0
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 0
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_141
timestamp 0
transform 1 0 14076 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_153
timestamp 0
transform 1 0 15180 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_165
timestamp 0
transform 1 0 16284 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_177
timestamp 0
transform 1 0 17388 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_189
timestamp 0
transform 1 0 18492 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 0
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 0
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_209
timestamp 0
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_221
timestamp 0
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_233
timestamp 0
transform 1 0 22540 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_245
timestamp 0
transform 1 0 23644 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_251
timestamp 0
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 0
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_265
timestamp 0
transform 1 0 25484 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_277
timestamp 0
transform 1 0 26588 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_289
timestamp 0
transform 1 0 27692 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_301
timestamp 0
transform 1 0 28796 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_307
timestamp 0
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_309
timestamp 0
transform 1 0 29532 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_321
timestamp 0
transform 1 0 30636 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_333
timestamp 0
transform 1 0 31740 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_345
timestamp 0
transform 1 0 32844 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_357
timestamp 0
transform 1 0 33948 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_363
timestamp 0
transform 1 0 34500 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_365
timestamp 0
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_377
timestamp 0
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_389
timestamp 0
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_401
timestamp 0
transform 1 0 37996 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 0
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 0
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_27
timestamp 0
transform 1 0 3588 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_39
timestamp 0
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_51
timestamp 0
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_55
timestamp 0
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_57
timestamp 0
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_69
timestamp 0
transform 1 0 7452 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_81
timestamp 0
transform 1 0 8556 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_93
timestamp 0
transform 1 0 9660 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_105
timestamp 0
transform 1 0 10764 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_111
timestamp 0
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_113
timestamp 0
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_125
timestamp 0
transform 1 0 12604 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_137
timestamp 0
transform 1 0 13708 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_149
timestamp 0
transform 1 0 14812 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_161
timestamp 0
transform 1 0 15916 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 0
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 0
transform 1 0 16652 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_181
timestamp 0
transform 1 0 17756 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_193
timestamp 0
transform 1 0 18860 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_205
timestamp 0
transform 1 0 19964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_217
timestamp 0
transform 1 0 21068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_223
timestamp 0
transform 1 0 21620 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_225
timestamp 0
transform 1 0 21804 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_237
timestamp 0
transform 1 0 22908 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_249
timestamp 0
transform 1 0 24012 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_261
timestamp 0
transform 1 0 25116 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_273
timestamp 0
transform 1 0 26220 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_279
timestamp 0
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 0
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 0
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_305
timestamp 0
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_317
timestamp 0
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_329
timestamp 0
transform 1 0 31372 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_335
timestamp 0
transform 1 0 31924 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_337
timestamp 0
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_349
timestamp 0
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_361
timestamp 0
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_373
timestamp 0
transform 1 0 35420 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_385
timestamp 0
transform 1 0 36524 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_391
timestamp 0
transform 1 0 37076 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_393
timestamp 0
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_405
timestamp 0
transform 1 0 38364 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 0
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 0
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 0
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_29
timestamp 0
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_41
timestamp 0
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_53
timestamp 0
transform 1 0 5980 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_65
timestamp 0
transform 1 0 7084 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_77
timestamp 0
transform 1 0 8188 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 0
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_85
timestamp 0
transform 1 0 8924 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_97
timestamp 0
transform 1 0 10028 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_109
timestamp 0
transform 1 0 11132 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_121
timestamp 0
transform 1 0 12236 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_133
timestamp 0
transform 1 0 13340 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 0
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 0
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_153
timestamp 0
transform 1 0 15180 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_165
timestamp 0
transform 1 0 16284 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_177
timestamp 0
transform 1 0 17388 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_189
timestamp 0
transform 1 0 18492 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_195
timestamp 0
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_197
timestamp 0
transform 1 0 19228 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_209
timestamp 0
transform 1 0 20332 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_221
timestamp 0
transform 1 0 21436 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_233
timestamp 0
transform 1 0 22540 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_245
timestamp 0
transform 1 0 23644 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_251
timestamp 0
transform 1 0 24196 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_253
timestamp 0
transform 1 0 24380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_265
timestamp 0
transform 1 0 25484 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_277
timestamp 0
transform 1 0 26588 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_289
timestamp 0
transform 1 0 27692 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_301
timestamp 0
transform 1 0 28796 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 0
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_309
timestamp 0
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_321
timestamp 0
transform 1 0 30636 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_333
timestamp 0
transform 1 0 31740 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_345
timestamp 0
transform 1 0 32844 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_357
timestamp 0
transform 1 0 33948 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_363
timestamp 0
transform 1 0 34500 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_365
timestamp 0
transform 1 0 34684 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_377
timestamp 0
transform 1 0 35788 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_389
timestamp 0
transform 1 0 36892 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_401
timestamp 0
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 0
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 0
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_27
timestamp 0
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_39
timestamp 0
transform 1 0 4692 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_51
timestamp 0
transform 1 0 5796 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 0
transform 1 0 6164 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 0
transform 1 0 6348 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_69
timestamp 0
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_81
timestamp 0
transform 1 0 8556 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_93
timestamp 0
transform 1 0 9660 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_105
timestamp 0
transform 1 0 10764 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_111
timestamp 0
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_113
timestamp 0
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_125
timestamp 0
transform 1 0 12604 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_137
timestamp 0
transform 1 0 13708 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_149
timestamp 0
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_161
timestamp 0
transform 1 0 15916 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 0
transform 1 0 16468 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_169
timestamp 0
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_181
timestamp 0
transform 1 0 17756 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_193
timestamp 0
transform 1 0 18860 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_205
timestamp 0
transform 1 0 19964 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_217
timestamp 0
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_223
timestamp 0
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_225
timestamp 0
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_237
timestamp 0
transform 1 0 22908 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_249
timestamp 0
transform 1 0 24012 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_261
timestamp 0
transform 1 0 25116 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_273
timestamp 0
transform 1 0 26220 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_279
timestamp 0
transform 1 0 26772 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_281
timestamp 0
transform 1 0 26956 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_293
timestamp 0
transform 1 0 28060 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_305
timestamp 0
transform 1 0 29164 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_317
timestamp 0
transform 1 0 30268 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_329
timestamp 0
transform 1 0 31372 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_335
timestamp 0
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_337
timestamp 0
transform 1 0 32108 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_349
timestamp 0
transform 1 0 33212 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_361
timestamp 0
transform 1 0 34316 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_373
timestamp 0
transform 1 0 35420 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_385
timestamp 0
transform 1 0 36524 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_391
timestamp 0
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_393
timestamp 0
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_405
timestamp 0
transform 1 0 38364 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 0
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 0
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 0
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_29
timestamp 0
transform 1 0 3772 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_41
timestamp 0
transform 1 0 4876 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_53
timestamp 0
transform 1 0 5980 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_65
timestamp 0
transform 1 0 7084 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_77
timestamp 0
transform 1 0 8188 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_83
timestamp 0
transform 1 0 8740 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_85
timestamp 0
transform 1 0 8924 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_97
timestamp 0
transform 1 0 10028 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_109
timestamp 0
transform 1 0 11132 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_121
timestamp 0
transform 1 0 12236 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_133
timestamp 0
transform 1 0 13340 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 0
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_141
timestamp 0
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_153
timestamp 0
transform 1 0 15180 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_165
timestamp 0
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_177
timestamp 0
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_189
timestamp 0
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_195
timestamp 0
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_197
timestamp 0
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_209
timestamp 0
transform 1 0 20332 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_221
timestamp 0
transform 1 0 21436 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_233
timestamp 0
transform 1 0 22540 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_245
timestamp 0
transform 1 0 23644 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_251
timestamp 0
transform 1 0 24196 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_253
timestamp 0
transform 1 0 24380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_265
timestamp 0
transform 1 0 25484 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_277
timestamp 0
transform 1 0 26588 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_289
timestamp 0
transform 1 0 27692 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_301
timestamp 0
transform 1 0 28796 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_307
timestamp 0
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_309
timestamp 0
transform 1 0 29532 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_321
timestamp 0
transform 1 0 30636 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_333
timestamp 0
transform 1 0 31740 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_345
timestamp 0
transform 1 0 32844 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_357
timestamp 0
transform 1 0 33948 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_363
timestamp 0
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_365
timestamp 0
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_377
timestamp 0
transform 1 0 35788 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_389
timestamp 0
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_401
timestamp 0
transform 1 0 37996 0 1 29376
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 0
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 0
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_27
timestamp 0
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_39
timestamp 0
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_51
timestamp 0
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 0
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_57
timestamp 0
transform 1 0 6348 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_69
timestamp 0
transform 1 0 7452 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_81
timestamp 0
transform 1 0 8556 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_93
timestamp 0
transform 1 0 9660 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_105
timestamp 0
transform 1 0 10764 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 0
transform 1 0 11316 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 0
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_125
timestamp 0
transform 1 0 12604 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_137
timestamp 0
transform 1 0 13708 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_149
timestamp 0
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_161
timestamp 0
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 0
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_169
timestamp 0
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_181
timestamp 0
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_193
timestamp 0
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_205
timestamp 0
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_217
timestamp 0
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_223
timestamp 0
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 0
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_237
timestamp 0
transform 1 0 22908 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_249
timestamp 0
transform 1 0 24012 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_261
timestamp 0
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_273
timestamp 0
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_279
timestamp 0
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 0
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_293
timestamp 0
transform 1 0 28060 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_305
timestamp 0
transform 1 0 29164 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_317
timestamp 0
transform 1 0 30268 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_329
timestamp 0
transform 1 0 31372 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_335
timestamp 0
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_337
timestamp 0
transform 1 0 32108 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_349
timestamp 0
transform 1 0 33212 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_361
timestamp 0
transform 1 0 34316 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_373
timestamp 0
transform 1 0 35420 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_385
timestamp 0
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_391
timestamp 0
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_393
timestamp 0
transform 1 0 37260 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_405
timestamp 0
transform 1 0 38364 0 -1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 0
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 0
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 0
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_29
timestamp 0
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_41
timestamp 0
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_53
timestamp 0
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_65
timestamp 0
transform 1 0 7084 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_77
timestamp 0
transform 1 0 8188 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_83
timestamp 0
transform 1 0 8740 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_85
timestamp 0
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_97
timestamp 0
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_109
timestamp 0
transform 1 0 11132 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_121
timestamp 0
transform 1 0 12236 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_133
timestamp 0
transform 1 0 13340 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_139
timestamp 0
transform 1 0 13892 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_141
timestamp 0
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_153
timestamp 0
transform 1 0 15180 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_165
timestamp 0
transform 1 0 16284 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_177
timestamp 0
transform 1 0 17388 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_189
timestamp 0
transform 1 0 18492 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_195
timestamp 0
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_197
timestamp 0
transform 1 0 19228 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_209
timestamp 0
transform 1 0 20332 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_221
timestamp 0
transform 1 0 21436 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_233
timestamp 0
transform 1 0 22540 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_245
timestamp 0
transform 1 0 23644 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_251
timestamp 0
transform 1 0 24196 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_253
timestamp 0
transform 1 0 24380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_265
timestamp 0
transform 1 0 25484 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_277
timestamp 0
transform 1 0 26588 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_289
timestamp 0
transform 1 0 27692 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_301
timestamp 0
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_307
timestamp 0
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_309
timestamp 0
transform 1 0 29532 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_321
timestamp 0
transform 1 0 30636 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_333
timestamp 0
transform 1 0 31740 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_345
timestamp 0
transform 1 0 32844 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_357
timestamp 0
transform 1 0 33948 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_363
timestamp 0
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_365
timestamp 0
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_377
timestamp 0
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_389
timestamp 0
transform 1 0 36892 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_401
timestamp 0
transform 1 0 37996 0 1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 0
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 0
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 0
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 0
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 0
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 0
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 0
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_69
timestamp 0
transform 1 0 7452 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_81
timestamp 0
transform 1 0 8556 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_93
timestamp 0
transform 1 0 9660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_105
timestamp 0
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_111
timestamp 0
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_113
timestamp 0
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_125
timestamp 0
transform 1 0 12604 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_137
timestamp 0
transform 1 0 13708 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_149
timestamp 0
transform 1 0 14812 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_161
timestamp 0
transform 1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_167
timestamp 0
transform 1 0 16468 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_169
timestamp 0
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_181
timestamp 0
transform 1 0 17756 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_193
timestamp 0
transform 1 0 18860 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_205
timestamp 0
transform 1 0 19964 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_217
timestamp 0
transform 1 0 21068 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_223
timestamp 0
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_225
timestamp 0
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_237
timestamp 0
transform 1 0 22908 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_249
timestamp 0
transform 1 0 24012 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_261
timestamp 0
transform 1 0 25116 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_273
timestamp 0
transform 1 0 26220 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 0
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_281
timestamp 0
transform 1 0 26956 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_293
timestamp 0
transform 1 0 28060 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_305
timestamp 0
transform 1 0 29164 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_317
timestamp 0
transform 1 0 30268 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_329
timestamp 0
transform 1 0 31372 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_335
timestamp 0
transform 1 0 31924 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_337
timestamp 0
transform 1 0 32108 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_349
timestamp 0
transform 1 0 33212 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_361
timestamp 0
transform 1 0 34316 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_373
timestamp 0
transform 1 0 35420 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_385
timestamp 0
transform 1 0 36524 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_391
timestamp 0
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_393
timestamp 0
transform 1 0 37260 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_405
timestamp 0
transform 1 0 38364 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 0
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 0
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 0
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_29
timestamp 0
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_41
timestamp 0
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_53
timestamp 0
transform 1 0 5980 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_65
timestamp 0
transform 1 0 7084 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_77
timestamp 0
transform 1 0 8188 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_83
timestamp 0
transform 1 0 8740 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 0
transform 1 0 8924 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_97
timestamp 0
transform 1 0 10028 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_109
timestamp 0
transform 1 0 11132 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_121
timestamp 0
transform 1 0 12236 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_133
timestamp 0
transform 1 0 13340 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_139
timestamp 0
transform 1 0 13892 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 0
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_153
timestamp 0
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_165
timestamp 0
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_177
timestamp 0
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_189
timestamp 0
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_195
timestamp 0
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_197
timestamp 0
transform 1 0 19228 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_209
timestamp 0
transform 1 0 20332 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_221
timestamp 0
transform 1 0 21436 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_233
timestamp 0
transform 1 0 22540 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_245
timestamp 0
transform 1 0 23644 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_251
timestamp 0
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_253
timestamp 0
transform 1 0 24380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_265
timestamp 0
transform 1 0 25484 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_277
timestamp 0
transform 1 0 26588 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_289
timestamp 0
transform 1 0 27692 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_301
timestamp 0
transform 1 0 28796 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_307
timestamp 0
transform 1 0 29348 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_309
timestamp 0
transform 1 0 29532 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_321
timestamp 0
transform 1 0 30636 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_333
timestamp 0
transform 1 0 31740 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_345
timestamp 0
transform 1 0 32844 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_357
timestamp 0
transform 1 0 33948 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_363
timestamp 0
transform 1 0 34500 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_365
timestamp 0
transform 1 0 34684 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_377
timestamp 0
transform 1 0 35788 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_389
timestamp 0
transform 1 0 36892 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_401
timestamp 0
transform 1 0 37996 0 1 31552
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 0
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 0
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 0
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_39
timestamp 0
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_51
timestamp 0
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_55
timestamp 0
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 0
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_69
timestamp 0
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_81
timestamp 0
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_93
timestamp 0
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_105
timestamp 0
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_111
timestamp 0
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_113
timestamp 0
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_125
timestamp 0
transform 1 0 12604 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_137
timestamp 0
transform 1 0 13708 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_149
timestamp 0
transform 1 0 14812 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_161
timestamp 0
transform 1 0 15916 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_167
timestamp 0
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_169
timestamp 0
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_181
timestamp 0
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_193
timestamp 0
transform 1 0 18860 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_205
timestamp 0
transform 1 0 19964 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_217
timestamp 0
transform 1 0 21068 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_223
timestamp 0
transform 1 0 21620 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_225
timestamp 0
transform 1 0 21804 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_237
timestamp 0
transform 1 0 22908 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_249
timestamp 0
transform 1 0 24012 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_261
timestamp 0
transform 1 0 25116 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_273
timestamp 0
transform 1 0 26220 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_279
timestamp 0
transform 1 0 26772 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_281
timestamp 0
transform 1 0 26956 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_293
timestamp 0
transform 1 0 28060 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_305
timestamp 0
transform 1 0 29164 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_317
timestamp 0
transform 1 0 30268 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_329
timestamp 0
transform 1 0 31372 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_335
timestamp 0
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_337
timestamp 0
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_349
timestamp 0
transform 1 0 33212 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_361
timestamp 0
transform 1 0 34316 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_373
timestamp 0
transform 1 0 35420 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_385
timestamp 0
transform 1 0 36524 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_391
timestamp 0
transform 1 0 37076 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_393
timestamp 0
transform 1 0 37260 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_405
timestamp 0
transform 1 0 38364 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 0
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 0
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 0
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_29
timestamp 0
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_41
timestamp 0
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_53
timestamp 0
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_65
timestamp 0
transform 1 0 7084 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_77
timestamp 0
transform 1 0 8188 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_83
timestamp 0
transform 1 0 8740 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_85
timestamp 0
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_97
timestamp 0
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_109
timestamp 0
transform 1 0 11132 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_121
timestamp 0
transform 1 0 12236 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_133
timestamp 0
transform 1 0 13340 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 0
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 0
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_153
timestamp 0
transform 1 0 15180 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_165
timestamp 0
transform 1 0 16284 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_177
timestamp 0
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_189
timestamp 0
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_195
timestamp 0
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_197
timestamp 0
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_209
timestamp 0
transform 1 0 20332 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_221
timestamp 0
transform 1 0 21436 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_233
timestamp 0
transform 1 0 22540 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_245
timestamp 0
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_251
timestamp 0
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_253
timestamp 0
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_265
timestamp 0
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_277
timestamp 0
transform 1 0 26588 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_289
timestamp 0
transform 1 0 27692 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_301
timestamp 0
transform 1 0 28796 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_307
timestamp 0
transform 1 0 29348 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_309
timestamp 0
transform 1 0 29532 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_321
timestamp 0
transform 1 0 30636 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_333
timestamp 0
transform 1 0 31740 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_345
timestamp 0
transform 1 0 32844 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_357
timestamp 0
transform 1 0 33948 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_363
timestamp 0
transform 1 0 34500 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_365
timestamp 0
transform 1 0 34684 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_377
timestamp 0
transform 1 0 35788 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_389
timestamp 0
transform 1 0 36892 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_401
timestamp 0
transform 1 0 37996 0 1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 0
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 0
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 0
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_39
timestamp 0
transform 1 0 4692 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_51
timestamp 0
transform 1 0 5796 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 0
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_57
timestamp 0
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_69
timestamp 0
transform 1 0 7452 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_81
timestamp 0
transform 1 0 8556 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_93
timestamp 0
transform 1 0 9660 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_105
timestamp 0
transform 1 0 10764 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 0
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 0
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 0
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_137
timestamp 0
transform 1 0 13708 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_149
timestamp 0
transform 1 0 14812 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_161
timestamp 0
transform 1 0 15916 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 0
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_169
timestamp 0
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_181
timestamp 0
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_193
timestamp 0
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_205
timestamp 0
transform 1 0 19964 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_217
timestamp 0
transform 1 0 21068 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_223
timestamp 0
transform 1 0 21620 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_225
timestamp 0
transform 1 0 21804 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_237
timestamp 0
transform 1 0 22908 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_249
timestamp 0
transform 1 0 24012 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_261
timestamp 0
transform 1 0 25116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_273
timestamp 0
transform 1 0 26220 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_279
timestamp 0
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_281
timestamp 0
transform 1 0 26956 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_293
timestamp 0
transform 1 0 28060 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_305
timestamp 0
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_317
timestamp 0
transform 1 0 30268 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_329
timestamp 0
transform 1 0 31372 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_335
timestamp 0
transform 1 0 31924 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_337
timestamp 0
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_349
timestamp 0
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_361
timestamp 0
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_373
timestamp 0
transform 1 0 35420 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_385
timestamp 0
transform 1 0 36524 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_391
timestamp 0
transform 1 0 37076 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_393
timestamp 0
transform 1 0 37260 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_401
timestamp 0
transform 1 0 37996 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 0
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 0
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 0
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_29
timestamp 0
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_41
timestamp 0
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_53
timestamp 0
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_65
timestamp 0
transform 1 0 7084 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_77
timestamp 0
transform 1 0 8188 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_83
timestamp 0
transform 1 0 8740 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_85
timestamp 0
transform 1 0 8924 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_97
timestamp 0
transform 1 0 10028 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_109
timestamp 0
transform 1 0 11132 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_121
timestamp 0
transform 1 0 12236 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_133
timestamp 0
transform 1 0 13340 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_139
timestamp 0
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_141
timestamp 0
transform 1 0 14076 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_153
timestamp 0
transform 1 0 15180 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_165
timestamp 0
transform 1 0 16284 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_177
timestamp 0
transform 1 0 17388 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_189
timestamp 0
transform 1 0 18492 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 0
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_197
timestamp 0
transform 1 0 19228 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_209
timestamp 0
transform 1 0 20332 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_221
timestamp 0
transform 1 0 21436 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_233
timestamp 0
transform 1 0 22540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_245
timestamp 0
transform 1 0 23644 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_251
timestamp 0
transform 1 0 24196 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_253
timestamp 0
transform 1 0 24380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_265
timestamp 0
transform 1 0 25484 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_277
timestamp 0
transform 1 0 26588 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_289
timestamp 0
transform 1 0 27692 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_301
timestamp 0
transform 1 0 28796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_307
timestamp 0
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_309
timestamp 0
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_321
timestamp 0
transform 1 0 30636 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_333
timestamp 0
transform 1 0 31740 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_345
timestamp 0
transform 1 0 32844 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_357
timestamp 0
transform 1 0 33948 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_363
timestamp 0
transform 1 0 34500 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_365
timestamp 0
transform 1 0 34684 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_377
timestamp 0
transform 1 0 35788 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_389
timestamp 0
transform 1 0 36892 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_401
timestamp 0
transform 1 0 37996 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 0
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 0
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 0
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_39
timestamp 0
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_51
timestamp 0
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 0
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 0
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_69
timestamp 0
transform 1 0 7452 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_81
timestamp 0
transform 1 0 8556 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_93
timestamp 0
transform 1 0 9660 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_105
timestamp 0
transform 1 0 10764 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 0
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_113
timestamp 0
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_125
timestamp 0
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_137
timestamp 0
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_149
timestamp 0
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_161
timestamp 0
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_167
timestamp 0
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_169
timestamp 0
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_181
timestamp 0
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_193
timestamp 0
transform 1 0 18860 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_205
timestamp 0
transform 1 0 19964 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_217
timestamp 0
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_223
timestamp 0
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_225
timestamp 0
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_237
timestamp 0
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_249
timestamp 0
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_261
timestamp 0
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_273
timestamp 0
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_279
timestamp 0
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_281
timestamp 0
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_293
timestamp 0
transform 1 0 28060 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_305
timestamp 0
transform 1 0 29164 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_317
timestamp 0
transform 1 0 30268 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_329
timestamp 0
transform 1 0 31372 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_335
timestamp 0
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_337
timestamp 0
transform 1 0 32108 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_349
timestamp 0
transform 1 0 33212 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_361
timestamp 0
transform 1 0 34316 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_373
timestamp 0
transform 1 0 35420 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_385
timestamp 0
transform 1 0 36524 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_391
timestamp 0
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_393
timestamp 0
transform 1 0 37260 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_405
timestamp 0
transform 1 0 38364 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_3
timestamp 0
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_15
timestamp 0
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 0
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 0
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 0
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_53
timestamp 0
transform 1 0 5980 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_65
timestamp 0
transform 1 0 7084 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_77
timestamp 0
transform 1 0 8188 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_83
timestamp 0
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_85
timestamp 0
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_97
timestamp 0
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_109
timestamp 0
transform 1 0 11132 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_121
timestamp 0
transform 1 0 12236 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_133
timestamp 0
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 0
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_141
timestamp 0
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_153
timestamp 0
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_165
timestamp 0
transform 1 0 16284 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_177
timestamp 0
transform 1 0 17388 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_189
timestamp 0
transform 1 0 18492 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_195
timestamp 0
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_197
timestamp 0
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_209
timestamp 0
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_221
timestamp 0
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_233
timestamp 0
transform 1 0 22540 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_245
timestamp 0
transform 1 0 23644 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_251
timestamp 0
transform 1 0 24196 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_253
timestamp 0
transform 1 0 24380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_265
timestamp 0
transform 1 0 25484 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_277
timestamp 0
transform 1 0 26588 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_289
timestamp 0
transform 1 0 27692 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_301
timestamp 0
transform 1 0 28796 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 0
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_309
timestamp 0
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_321
timestamp 0
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_333
timestamp 0
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_345
timestamp 0
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_357
timestamp 0
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_363
timestamp 0
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_365
timestamp 0
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_377
timestamp 0
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_389
timestamp 0
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_401
timestamp 0
transform 1 0 37996 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 0
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 0
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 0
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_39
timestamp 0
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 0
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 0
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_57
timestamp 0
transform 1 0 6348 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_69
timestamp 0
transform 1 0 7452 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_81
timestamp 0
transform 1 0 8556 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_93
timestamp 0
transform 1 0 9660 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_105
timestamp 0
transform 1 0 10764 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_111
timestamp 0
transform 1 0 11316 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 0
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_125
timestamp 0
transform 1 0 12604 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_137
timestamp 0
transform 1 0 13708 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_149
timestamp 0
transform 1 0 14812 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_161
timestamp 0
transform 1 0 15916 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_167
timestamp 0
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_169
timestamp 0
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_181
timestamp 0
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_193
timestamp 0
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_205
timestamp 0
transform 1 0 19964 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_217
timestamp 0
transform 1 0 21068 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 0
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_225
timestamp 0
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_237
timestamp 0
transform 1 0 22908 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_249
timestamp 0
transform 1 0 24012 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_261
timestamp 0
transform 1 0 25116 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_273
timestamp 0
transform 1 0 26220 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_279
timestamp 0
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_281
timestamp 0
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_293
timestamp 0
transform 1 0 28060 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_305
timestamp 0
transform 1 0 29164 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_317
timestamp 0
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_329
timestamp 0
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_335
timestamp 0
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_337
timestamp 0
transform 1 0 32108 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_349
timestamp 0
transform 1 0 33212 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_361
timestamp 0
transform 1 0 34316 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_373
timestamp 0
transform 1 0 35420 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_385
timestamp 0
transform 1 0 36524 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_391
timestamp 0
transform 1 0 37076 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_393
timestamp 0
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_405
timestamp 0
transform 1 0 38364 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_3
timestamp 0
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_15
timestamp 0
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 0
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 0
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_41
timestamp 0
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_53
timestamp 0
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_65
timestamp 0
transform 1 0 7084 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_77
timestamp 0
transform 1 0 8188 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_83
timestamp 0
transform 1 0 8740 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_85
timestamp 0
transform 1 0 8924 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_97
timestamp 0
transform 1 0 10028 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_109
timestamp 0
transform 1 0 11132 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_121
timestamp 0
transform 1 0 12236 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_133
timestamp 0
transform 1 0 13340 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_139
timestamp 0
transform 1 0 13892 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_141
timestamp 0
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_153
timestamp 0
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_165
timestamp 0
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_177
timestamp 0
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_189
timestamp 0
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_195
timestamp 0
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_197
timestamp 0
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_209
timestamp 0
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_221
timestamp 0
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_233
timestamp 0
transform 1 0 22540 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_245
timestamp 0
transform 1 0 23644 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_251
timestamp 0
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_253
timestamp 0
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_265
timestamp 0
transform 1 0 25484 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_277
timestamp 0
transform 1 0 26588 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_289
timestamp 0
transform 1 0 27692 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_301
timestamp 0
transform 1 0 28796 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_307
timestamp 0
transform 1 0 29348 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_309
timestamp 0
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_321
timestamp 0
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_333
timestamp 0
transform 1 0 31740 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_345
timestamp 0
transform 1 0 32844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_357
timestamp 0
transform 1 0 33948 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_363
timestamp 0
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_365
timestamp 0
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_377
timestamp 0
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_389
timestamp 0
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_401
timestamp 0
transform 1 0 37996 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 0
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 0
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 0
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 0
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 0
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 0
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_57
timestamp 0
transform 1 0 6348 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_69
timestamp 0
transform 1 0 7452 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_81
timestamp 0
transform 1 0 8556 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_93
timestamp 0
transform 1 0 9660 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_105
timestamp 0
transform 1 0 10764 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_111
timestamp 0
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_113
timestamp 0
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_125
timestamp 0
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_137
timestamp 0
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_149
timestamp 0
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_161
timestamp 0
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_167
timestamp 0
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_169
timestamp 0
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_181
timestamp 0
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_193
timestamp 0
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_205
timestamp 0
transform 1 0 19964 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_217
timestamp 0
transform 1 0 21068 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_223
timestamp 0
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_225
timestamp 0
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_237
timestamp 0
transform 1 0 22908 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_249
timestamp 0
transform 1 0 24012 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_261
timestamp 0
transform 1 0 25116 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_273
timestamp 0
transform 1 0 26220 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_279
timestamp 0
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_281
timestamp 0
transform 1 0 26956 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_293
timestamp 0
transform 1 0 28060 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_305
timestamp 0
transform 1 0 29164 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_317
timestamp 0
transform 1 0 30268 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_329
timestamp 0
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_335
timestamp 0
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_337
timestamp 0
transform 1 0 32108 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_349
timestamp 0
transform 1 0 33212 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_361
timestamp 0
transform 1 0 34316 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_373
timestamp 0
transform 1 0 35420 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_385
timestamp 0
transform 1 0 36524 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_391
timestamp 0
transform 1 0 37076 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_393
timestamp 0
transform 1 0 37260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_405
timestamp 0
transform 1 0 38364 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_9
timestamp 0
transform 1 0 1932 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_21
timestamp 0
transform 1 0 3036 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 0
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 0
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 0
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_53
timestamp 0
transform 1 0 5980 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_57
timestamp 0
transform 1 0 6348 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_69
timestamp 0
transform 1 0 7452 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_81
timestamp 0
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_85
timestamp 0
transform 1 0 8924 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_93
timestamp 0
transform 1 0 9660 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_100
timestamp 0
transform 1 0 10304 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_113
timestamp 0
transform 1 0 11500 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_125
timestamp 0
transform 1 0 12604 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_137
timestamp 0
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_141
timestamp 0
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_153
timestamp 0
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_165
timestamp 0
transform 1 0 16284 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_169
timestamp 0
transform 1 0 16652 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_181
timestamp 0
transform 1 0 17756 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_193
timestamp 0
transform 1 0 18860 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_197
timestamp 0
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_209
timestamp 0
transform 1 0 20332 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_221
timestamp 0
transform 1 0 21436 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_225
timestamp 0
transform 1 0 21804 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_237
timestamp 0
transform 1 0 22908 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_249
timestamp 0
transform 1 0 24012 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_253
timestamp 0
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_265
timestamp 0
transform 1 0 25484 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_277
timestamp 0
transform 1 0 26588 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_281
timestamp 0
transform 1 0 26956 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_293
timestamp 0
transform 1 0 28060 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_305
timestamp 0
transform 1 0 29164 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_309
timestamp 0
transform 1 0 29532 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_321
timestamp 0
transform 1 0 30636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_333
timestamp 0
transform 1 0 31740 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_337
timestamp 0
transform 1 0 32108 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_349
timestamp 0
transform 1 0 33212 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_357
timestamp 0
transform 1 0 33948 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_363
timestamp 0
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_365
timestamp 0
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_377
timestamp 0
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_389
timestamp 0
transform 1 0 36892 0 1 36992
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_393
timestamp 0
transform 1 0 37260 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_405
timestamp 0
transform 1 0 38364 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1
timestamp 0
transform -1 0 25576 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 0
transform -1 0 30268 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 0
transform 1 0 30268 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 0
transform 1 0 26220 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 0
transform -1 0 27692 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 0
transform -1 0 28888 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 0
transform -1 0 27692 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 0
transform -1 0 22816 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 0
transform 1 0 23460 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 0
transform -1 0 27876 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 0
transform 1 0 22540 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 0
transform 1 0 23184 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 0
transform -1 0 23552 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 0
transform 1 0 23552 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold15
timestamp 0
transform 1 0 28336 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold16
timestamp 0
transform -1 0 23460 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold17
timestamp 0
transform -1 0 24288 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold18
timestamp 0
transform -1 0 25116 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold19
timestamp 0
transform -1 0 23092 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold20
timestamp 0
transform -1 0 21160 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold21
timestamp 0
transform -1 0 24840 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold22
timestamp 0
transform -1 0 23000 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold23
timestamp 0
transform -1 0 23184 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold24
timestamp 0
transform -1 0 27692 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold25
timestamp 0
transform -1 0 20332 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold26
timestamp 0
transform -1 0 21160 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  input1
timestamp 0
transform -1 0 24196 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 0
transform -1 0 33948 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 0
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 0
transform 1 0 1380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 0
transform -1 0 35880 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 0
transform 1 0 1380 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input7
timestamp 0
transform 1 0 21988 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input8
timestamp 0
transform -1 0 38548 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 0
transform 1 0 11684 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 0
transform -1 0 38548 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output11
timestamp 0
transform -1 0 1932 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output12
timestamp 0
transform -1 0 10304 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 0
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 0
transform -1 0 38824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 0
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 0
transform -1 0 38824 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 0
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 0
transform -1 0 38824 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 0
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 0
transform -1 0 38824 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 0
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 0
transform -1 0 38824 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 0
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 0
transform -1 0 38824 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 0
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 0
transform -1 0 38824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 0
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 0
transform -1 0 38824 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 0
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 0
transform -1 0 38824 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 0
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 0
transform -1 0 38824 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 0
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 0
transform -1 0 38824 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 0
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 0
transform -1 0 38824 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 0
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 0
transform -1 0 38824 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 0
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 0
transform -1 0 38824 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 0
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 0
transform -1 0 38824 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 0
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 0
transform -1 0 38824 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 0
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 0
transform -1 0 38824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 0
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 0
transform -1 0 38824 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 0
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 0
transform -1 0 38824 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 0
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 0
transform -1 0 38824 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 0
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 0
transform -1 0 38824 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 0
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 0
transform -1 0 38824 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 0
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 0
transform -1 0 38824 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 0
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 0
transform -1 0 38824 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 0
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 0
transform -1 0 38824 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 0
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 0
transform -1 0 38824 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 0
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 0
transform -1 0 38824 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 0
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 0
transform -1 0 38824 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 0
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 0
transform -1 0 38824 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 0
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 0
transform -1 0 38824 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 0
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 0
transform -1 0 38824 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 0
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 0
transform -1 0 38824 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 0
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 0
transform -1 0 38824 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 0
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 0
transform -1 0 38824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 0
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 0
transform -1 0 38824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 0
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 0
transform -1 0 38824 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 0
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 0
transform -1 0 38824 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 0
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 0
transform -1 0 38824 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 0
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 0
transform -1 0 38824 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 0
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 0
transform -1 0 38824 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 0
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 0
transform -1 0 38824 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 0
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 0
transform -1 0 38824 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 0
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 0
transform -1 0 38824 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 0
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 0
transform -1 0 38824 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 0
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 0
transform -1 0 38824 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 0
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 0
transform -1 0 38824 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 0
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 0
transform -1 0 38824 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 0
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 0
transform -1 0 38824 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 0
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 0
transform -1 0 38824 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 0
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 0
transform -1 0 38824 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 0
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 0
transform -1 0 38824 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 0
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 0
transform -1 0 38824 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 0
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 0
transform -1 0 38824 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 0
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 0
transform -1 0 38824 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 0
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 0
transform -1 0 38824 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 0
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 0
transform -1 0 38824 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 0
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 0
transform -1 0 38824 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 0
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 0
transform -1 0 38824 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 0
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 0
transform -1 0 38824 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 0
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 0
transform -1 0 38824 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 0
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 0
transform -1 0 38824 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 0
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 0
transform -1 0 38824 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 0
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 0
transform -1 0 38824 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 0
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 0
transform -1 0 38824 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 0
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 0
transform -1 0 38824 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 0
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 0
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 0
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 0
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 0
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 0
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 0
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 0
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 0
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 0
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 0
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 0
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 0
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 0
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 0
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 0
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 0
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 0
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 0
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 0
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 0
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 0
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 0
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 0
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 0
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 0
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 0
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 0
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 0
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 0
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 0
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 0
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 0
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 0
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 0
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 0
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 0
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 0
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 0
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 0
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 0
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 0
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 0
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 0
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 0
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 0
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 0
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 0
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 0
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 0
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 0
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 0
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 0
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 0
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 0
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 0
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 0
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 0
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 0
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 0
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 0
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 0
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 0
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 0
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 0
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 0
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 0
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 0
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 0
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 0
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 0
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 0
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 0
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 0
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 0
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 0
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 0
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 0
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 0
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 0
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 0
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 0
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 0
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 0
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 0
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 0
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 0
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 0
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 0
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 0
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 0
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 0
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 0
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 0
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 0
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 0
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 0
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 0
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 0
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 0
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 0
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 0
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 0
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 0
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 0
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 0
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 0
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 0
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 0
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 0
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 0
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 0
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 0
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 0
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 0
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 0
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 0
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 0
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 0
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 0
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 0
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 0
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 0
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 0
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 0
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 0
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 0
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 0
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 0
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 0
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 0
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 0
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 0
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 0
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 0
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 0
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 0
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 0
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 0
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 0
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 0
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 0
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 0
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 0
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 0
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 0
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 0
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 0
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 0
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 0
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 0
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 0
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 0
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 0
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 0
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 0
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 0
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 0
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 0
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 0
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 0
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 0
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 0
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 0
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 0
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 0
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 0
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 0
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 0
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 0
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 0
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 0
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 0
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 0
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 0
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 0
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 0
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 0
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 0
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 0
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 0
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 0
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 0
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 0
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 0
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 0
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 0
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 0
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 0
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 0
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 0
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 0
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 0
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 0
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 0
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 0
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 0
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 0
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 0
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 0
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 0
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 0
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 0
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 0
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 0
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 0
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 0
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 0
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 0
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 0
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 0
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 0
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 0
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 0
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 0
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 0
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 0
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 0
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 0
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 0
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 0
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 0
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 0
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 0
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 0
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 0
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 0
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 0
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 0
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 0
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 0
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 0
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 0
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 0
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 0
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 0
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 0
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 0
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 0
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 0
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 0
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 0
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 0
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 0
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 0
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 0
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 0
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 0
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 0
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 0
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 0
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 0
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 0
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 0
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 0
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 0
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 0
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 0
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 0
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 0
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 0
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 0
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 0
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 0
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 0
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 0
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 0
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 0
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 0
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 0
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 0
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 0
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 0
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 0
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 0
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 0
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 0
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 0
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 0
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 0
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 0
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 0
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 0
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 0
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 0
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 0
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 0
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 0
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 0
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 0
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 0
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 0
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 0
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 0
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 0
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 0
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 0
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 0
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 0
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 0
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 0
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 0
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 0
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 0
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 0
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 0
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 0
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 0
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 0
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 0
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 0
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 0
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 0
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 0
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 0
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 0
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 0
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 0
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 0
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 0
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 0
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 0
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 0
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 0
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 0
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 0
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 0
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 0
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 0
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 0
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 0
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 0
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 0
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 0
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 0
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 0
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 0
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 0
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 0
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 0
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 0
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 0
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 0
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 0
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 0
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 0
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 0
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 0
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 0
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 0
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 0
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 0
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 0
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 0
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 0
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 0
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 0
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 0
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 0
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 0
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 0
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 0
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 0
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 0
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 0
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 0
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 0
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 0
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 0
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 0
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 0
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 0
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 0
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 0
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 0
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 0
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 0
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 0
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 0
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 0
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 0
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 0
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 0
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 0
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 0
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 0
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 0
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 0
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 0
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 0
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 0
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 0
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 0
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 0
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 0
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 0
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 0
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 0
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 0
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 0
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 0
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 0
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 0
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 0
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 0
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 0
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 0
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 0
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 0
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 0
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 0
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 0
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 0
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 0
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 0
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 0
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 0
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 0
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 0
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 0
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 0
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 0
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 0
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 0
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 0
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 0
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 0
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 0
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 0
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 0
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 0
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 0
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 0
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 0
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 0
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 0
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 0
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 0
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 0
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 0
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 0
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 0
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 0
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 0
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 0
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 0
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 0
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 0
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 0
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 0
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 0
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 0
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 0
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 0
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 0
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 0
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 0
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 0
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 0
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 0
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 0
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 0
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 0
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 0
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 0
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 0
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 0
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 0
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 0
transform 1 0 37168 0 1 36992
box -38 -48 130 592
<< labels >>
rlabel metal1 s 19964 36992 19964 36992 4 VGND
rlabel metal1 s 19964 37536 19964 37536 4 VPWR
rlabel metal1 s 25162 14008 25162 14008 4 _000_
rlabel metal1 s 25300 13294 25300 13294 4 _001_
rlabel metal2 s 27922 14178 27922 14178 4 _002_
rlabel metal1 s 27876 12410 27876 12410 4 _003_
rlabel metal1 s 28014 10710 28014 10710 4 _004_
rlabel metal2 s 27830 11492 27830 11492 4 _005_
rlabel metal1 s 24196 6358 24196 6358 4 _006_
rlabel metal1 s 26588 5338 26588 5338 4 _007_
rlabel metal1 s 25208 5746 25208 5746 4 _008_
rlabel metal1 s 29164 6222 29164 6222 4 _009_
rlabel metal1 s 29348 7310 29348 7310 4 _010_
rlabel metal1 s 29946 8058 29946 8058 4 _011_
rlabel metal1 s 25208 8398 25208 8398 4 _012_
rlabel metal1 s 26082 8874 26082 8874 4 _013_
rlabel metal2 s 27738 9758 27738 9758 4 _014_
rlabel metal2 s 21482 8738 21482 8738 4 _015_
rlabel metal1 s 24242 9146 24242 9146 4 _016_
rlabel metal1 s 21298 6630 21298 6630 4 _017_
rlabel metal1 s 22356 5338 22356 5338 4 _018_
rlabel metal2 s 23690 6188 23690 6188 4 _019_
rlabel metal1 s 20509 6970 20509 6970 4 _020_
rlabel metal1 s 22402 8058 22402 8058 4 _021_
rlabel metal1 s 21160 10778 21160 10778 4 _022_
rlabel metal1 s 22126 10744 22126 10744 4 _023_
rlabel metal2 s 23782 11220 23782 11220 4 _024_
rlabel metal2 s 23230 13668 23230 13668 4 _025_
rlabel metal1 s 22816 14450 22816 14450 4 _026_
rlabel metal1 s 18860 13974 18860 13974 4 _027_
rlabel metal1 s 18630 11662 18630 11662 4 _028_
rlabel metal1 s 21252 12954 21252 12954 4 _029_
rlabel metal1 s 19458 12614 19458 12614 4 _030_
rlabel metal1 s 20378 15062 20378 15062 4 _031_
rlabel metal1 s 21068 14314 21068 14314 4 _032_
rlabel metal1 s 28750 6868 28750 6868 4 _033_
rlabel metal1 s 25990 9554 25990 9554 4 _034_
rlabel metal1 s 23506 7514 23506 7514 4 _035_
rlabel metal1 s 25484 10030 25484 10030 4 _036_
rlabel metal1 s 29486 9962 29486 9962 4 _037_
rlabel metal1 s 26818 9588 26818 9588 4 _038_
rlabel metal1 s 26128 10642 26128 10642 4 _039_
rlabel metal1 s 25162 12614 25162 12614 4 _040_
rlabel metal1 s 25852 9622 25852 9622 4 _041_
rlabel metal2 s 27370 10880 27370 10880 4 _042_
rlabel metal2 s 26450 10880 26450 10880 4 _043_
rlabel metal1 s 27508 11866 27508 11866 4 _044_
rlabel metal1 s 30038 6732 30038 6732 4 _045_
rlabel metal1 s 27784 11186 27784 11186 4 _046_
rlabel metal1 s 27738 10778 27738 10778 4 _047_
rlabel metal1 s 25392 11526 25392 11526 4 _048_
rlabel metal1 s 26910 9350 26910 9350 4 _049_
rlabel metal1 s 23460 9690 23460 9690 4 _050_
rlabel metal2 s 24886 7174 24886 7174 4 _051_
rlabel metal1 s 26864 4794 26864 4794 4 _052_
rlabel metal1 s 26128 5338 26128 5338 4 _053_
rlabel metal1 s 26220 6698 26220 6698 4 _054_
rlabel metal1 s 29210 5644 29210 5644 4 _055_
rlabel metal1 s 28842 5338 28842 5338 4 _056_
rlabel metal1 s 28106 7888 28106 7888 4 _057_
rlabel metal1 s 28934 5712 28934 5712 4 _058_
rlabel metal1 s 28474 7276 28474 7276 4 _059_
rlabel metal1 s 29302 7514 29302 7514 4 _060_
rlabel metal2 s 30038 7412 30038 7412 4 _061_
rlabel metal2 s 29578 8364 29578 8364 4 _062_
rlabel metal1 s 27600 7242 27600 7242 4 _063_
rlabel metal1 s 26174 8432 26174 8432 4 _064_
rlabel metal1 s 29072 9010 29072 9010 4 _065_
rlabel metal1 s 28474 9962 28474 9962 4 _066_
rlabel metal1 s 27508 9010 27508 9010 4 _067_
rlabel metal1 s 21712 8466 21712 8466 4 _068_
rlabel metal1 s 24334 8942 24334 8942 4 _069_
rlabel metal1 s 21804 7378 21804 7378 4 _070_
rlabel metal1 s 23552 5202 23552 5202 4 _071_
rlabel metal1 s 23736 6766 23736 6766 4 _072_
rlabel metal1 s 20746 7412 20746 7412 4 _073_
rlabel metal1 s 22862 7922 22862 7922 4 _074_
rlabel metal1 s 25208 9350 25208 9350 4 _075_
rlabel metal2 s 25162 11458 25162 11458 4 _076_
rlabel metal1 s 24472 10506 24472 10506 4 _077_
rlabel metal1 s 21666 10642 21666 10642 4 _078_
rlabel metal2 s 23230 11067 23230 11067 4 _079_
rlabel metal2 s 23506 10608 23506 10608 4 _080_
rlabel metal2 s 25714 10132 25714 10132 4 _081_
rlabel metal2 s 23966 10812 23966 10812 4 _082_
rlabel metal1 s 23460 13294 23460 13294 4 _083_
rlabel metal1 s 23230 14994 23230 14994 4 _084_
rlabel metal1 s 19136 14586 19136 14586 4 _085_
rlabel metal1 s 18216 12206 18216 12206 4 _086_
rlabel metal1 s 21528 12410 21528 12410 4 _087_
rlabel metal1 s 19320 12818 19320 12818 4 _088_
rlabel metal1 s 21482 15130 21482 15130 4 _089_
rlabel metal1 s 21528 15470 21528 15470 4 _090_
rlabel metal1 s 24610 15538 24610 15538 4 _091_
rlabel metal1 s 24150 15538 24150 15538 4 _092_
rlabel metal1 s 25024 14994 25024 14994 4 _093_
rlabel metal1 s 20884 13430 20884 13430 4 _094_
rlabel metal1 s 20838 13498 20838 13498 4 _095_
rlabel metal1 s 23414 13702 23414 13702 4 _096_
rlabel metal1 s 25530 14382 25530 14382 4 _097_
rlabel metal1 s 29026 11220 29026 11220 4 _098_
rlabel metal2 s 28106 12274 28106 12274 4 _099_
rlabel metal1 s 19504 12410 19504 12410 4 _100_
rlabel metal1 s 25392 14246 25392 14246 4 _101_
rlabel metal1 s 27002 11662 27002 11662 4 _102_
rlabel metal2 s 23782 12517 23782 12517 4 _103_
rlabel metal1 s 25622 12240 25622 12240 4 _104_
rlabel metal1 s 24150 12410 24150 12410 4 _105_
rlabel metal1 s 25254 12138 25254 12138 4 _106_
rlabel metal1 s 25898 12852 25898 12852 4 _107_
rlabel metal1 s 26726 11798 26726 11798 4 _108_
rlabel metal1 s 25438 11186 25438 11186 4 _109_
rlabel metal1 s 25944 11186 25944 11186 4 _110_
rlabel metal1 s 27646 13498 27646 13498 4 _111_
rlabel metal1 s 24886 11118 24886 11118 4 bit_idx\[0\]
rlabel metal1 s 22862 11764 22862 11764 4 bit_idx\[1\]
rlabel metal1 s 24702 11526 24702 11526 4 bit_idx\[2\]
rlabel metal3 s 37567 21148 37567 21148 4 clk
rlabel metal1 s 27324 6630 27324 6630 4 clk_cnt\[0\]
rlabel metal2 s 23046 9010 23046 9010 4 clk_cnt\[10\]
rlabel metal1 s 23276 7310 23276 7310 4 clk_cnt\[11\]
rlabel metal2 s 23690 7072 23690 7072 4 clk_cnt\[12\]
rlabel metal1 s 22782 6766 22782 6766 4 clk_cnt\[13\]
rlabel metal1 s 22862 7310 22862 7310 4 clk_cnt\[14\]
rlabel metal2 s 23598 8092 23598 8092 4 clk_cnt\[15\]
rlabel metal1 s 27416 6766 27416 6766 4 clk_cnt\[1\]
rlabel metal2 s 26634 6324 26634 6324 4 clk_cnt\[2\]
rlabel metal1 s 28842 6698 28842 6698 4 clk_cnt\[3\]
rlabel metal2 s 30314 7684 30314 7684 4 clk_cnt\[4\]
rlabel metal1 s 28014 7242 28014 7242 4 clk_cnt\[5\]
rlabel metal1 s 27646 8500 27646 8500 4 clk_cnt\[6\]
rlabel metal1 s 26358 8874 26358 8874 4 clk_cnt\[7\]
rlabel metal1 s 29670 9690 29670 9690 4 clk_cnt\[8\]
rlabel metal1 s 23138 9146 23138 9146 4 clk_cnt\[9\]
rlabel metal1 s 22540 9962 22540 9962 4 clknet_0_clk
rlabel metal1 s 21942 6154 21942 6154 4 clknet_2_0__leaf_clk
rlabel metal1 s 18676 11730 18676 11730 4 clknet_2_1__leaf_clk
rlabel metal1 s 27738 10574 27738 10574 4 clknet_2_2__leaf_clk
rlabel metal2 s 27554 10948 27554 10948 4 clknet_2_3__leaf_clk
rlabel metal2 s 23874 1588 23874 1588 4 data_in[0]
rlabel metal1 s 33672 37230 33672 37230 4 data_in[1]
rlabel metal3 s 820 25228 820 25228 4 data_in[2]
rlabel metal2 s 46 1554 46 1554 4 data_in[3]
rlabel metal2 s 35466 1520 35466 1520 4 data_in[4]
rlabel metal3 s 1050 12308 1050 12308 4 data_in[5]
rlabel metal1 s 21988 37298 21988 37298 4 data_in[6]
rlabel metal1 s 38640 33490 38640 33490 4 data_in[7]
rlabel metal1 s 24978 13702 24978 13702 4 data_reg\[0\]
rlabel metal1 s 24656 14518 24656 14518 4 data_reg\[1\]
rlabel metal2 s 22218 13328 22218 13328 4 data_reg\[2\]
rlabel metal3 s 20470 11883 20470 11883 4 data_reg\[3\]
rlabel metal1 s 22816 13158 22816 13158 4 data_reg\[4\]
rlabel metal1 s 21068 12410 21068 12410 4 data_reg\[5\]
rlabel metal1 s 23000 15470 23000 15470 4 data_reg\[6\]
rlabel metal2 s 22402 15300 22402 15300 4 data_reg\[7\]
rlabel metal1 s 24104 2618 24104 2618 4 net1
rlabel metal1 s 38272 8602 38272 8602 4 net10
rlabel metal1 s 4347 37162 4347 37162 4 net11
rlabel metal1 s 23046 13260 23046 13260 4 net12
rlabel metal1 s 22179 14314 22179 14314 4 net13
rlabel metal1 s 23085 9622 23085 9622 4 net14
rlabel metal1 s 26549 13974 26549 13974 4 net15
rlabel metal2 s 26266 12852 26266 12852 4 net16
rlabel metal1 s 24058 10676 24058 10676 4 net17
rlabel metal1 s 29279 10030 29279 10030 4 net18
rlabel metal1 s 30774 8058 30774 8058 4 net19
rlabel metal2 s 23690 15606 23690 15606 4 net2
rlabel metal1 s 27094 9010 27094 9010 4 net20
rlabel metal1 s 26680 6426 26680 6426 4 net21
rlabel metal1 s 28336 5202 28336 5202 4 net22
rlabel metal1 s 26818 8398 26818 8398 4 net23
rlabel metal1 s 21896 7310 21896 7310 4 net24
rlabel metal1 s 24104 8058 24104 8058 4 net25
rlabel metal1 s 26772 5202 26772 5202 4 net26
rlabel metal1 s 23828 6698 23828 6698 4 net27
rlabel metal1 s 24242 9078 24242 9078 4 net28
rlabel metal1 s 20838 7276 20838 7276 4 net29
rlabel metal1 s 4301 25194 4301 25194 4 net3
rlabel metal1 s 24518 6834 24518 6834 4 net30
rlabel metal1 s 29486 7854 29486 7854 4 net31
rlabel metal1 s 22632 9554 22632 9554 4 net32
rlabel metal1 s 23552 11118 23552 11118 4 net33
rlabel metal1 s 24196 13294 24196 13294 4 net34
rlabel metal1 s 22218 12070 22218 12070 4 net35
rlabel metal1 s 20194 12818 20194 12818 4 net36
rlabel metal1 s 23966 14994 23966 14994 4 net37
rlabel metal1 s 22126 15572 22126 15572 4 net38
rlabel metal1 s 22402 15130 22402 15130 4 net39
rlabel metal1 s 19090 12138 19090 12138 4 net4
rlabel metal2 s 25806 14144 25806 14144 4 net40
rlabel metal1 s 19228 11322 19228 11322 4 net41
rlabel metal1 s 20102 14042 20102 14042 4 net42
rlabel metal1 s 21988 12206 21988 12206 4 net5
rlabel metal1 s 4255 12614 4255 12614 4 net6
rlabel metal1 s 22816 15538 22816 15538 4 net7
rlabel metal1 s 23414 15436 23414 15436 4 net8
rlabel metal1 s 25806 12682 25806 12682 4 net9
rlabel metal1 s 27094 13838 27094 13838 4 parity_bit
rlabel metal2 s 11638 959 11638 959 4 rst_n
rlabel metal1 s 29532 12750 29532 12750 4 state\[0\]
rlabel metal2 s 29670 10948 29670 10948 4 state\[1\]
rlabel metal2 s 26818 12619 26818 12619 4 state\[2\]
rlabel metal3 s 820 37468 820 37468 4 tx_busy
rlabel metal1 s 9798 37434 9798 37434 4 tx_out
rlabel metal1 s 38640 8466 38640 8466 4 tx_start
flabel metal5 s 1056 36642 38872 36962 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal5 s 1056 6006 38872 6326 0 FreeSans 3200 0 0 0 VGND
port 1 nsew
flabel metal4 s 35588 2128 35908 37584 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal4 s 4868 2128 5188 37584 0 FreeSans 2400 90 0 0 VGND
port 1 nsew
flabel metal5 s 1056 35982 38872 36302 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal5 s 1056 5346 38872 5666 0 FreeSans 3200 0 0 0 VPWR
port 2 nsew
flabel metal4 s 34928 2128 35248 37584 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal4 s 4208 2128 4528 37584 0 FreeSans 2400 90 0 0 VPWR
port 2 nsew
flabel metal3 s 39200 21088 40000 21208 0 FreeSans 600 0 0 0 clk
port 3 nsew
flabel metal2 s 23846 0 23902 800 0 FreeSans 280 90 0 0 data_in[0]
port 4 nsew
flabel metal2 s 33506 39200 33562 40000 0 FreeSans 280 90 0 0 data_in[1]
port 5 nsew
flabel metal3 s 0 25168 800 25288 0 FreeSans 600 0 0 0 data_in[2]
port 6 nsew
flabel metal2 s 18 0 74 800 0 FreeSans 280 90 0 0 data_in[3]
port 7 nsew
flabel metal2 s 35438 0 35494 800 0 FreeSans 280 90 0 0 data_in[4]
port 8 nsew
flabel metal3 s 0 12248 800 12368 0 FreeSans 600 0 0 0 data_in[5]
port 9 nsew
flabel metal2 s 21914 39200 21970 40000 0 FreeSans 280 90 0 0 data_in[6]
port 10 nsew
flabel metal3 s 39200 33328 40000 33448 0 FreeSans 600 0 0 0 data_in[7]
port 11 nsew
flabel metal2 s 11610 0 11666 800 0 FreeSans 280 90 0 0 rst_n
port 12 nsew
flabel metal3 s 0 37408 800 37528 0 FreeSans 600 0 0 0 tx_busy
port 13 nsew
flabel metal2 s 9678 39200 9734 40000 0 FreeSans 280 90 0 0 tx_out
port 14 nsew
flabel metal3 s 39200 8168 40000 8288 0 FreeSans 600 0 0 0 tx_start
port 15 nsew
<< properties >>
string FIXED_BBOX 0 0 40000 40000
<< end >>
