magic
tech sky130A
magscale 1 2
timestamp 1765484839
<< obsli1 >>
rect 1104 2159 38824 37553
<< obsm1 >>
rect 14 2128 38902 37584
<< metal2 >>
rect 9678 39200 9734 40000
rect 21914 39200 21970 40000
rect 33506 39200 33562 40000
rect 18 0 74 800
rect 11610 0 11666 800
rect 23846 0 23902 800
rect 35438 0 35494 800
<< obsm2 >>
rect 20 39144 9622 39200
rect 9790 39144 21858 39200
rect 22026 39144 33450 39200
rect 33618 39144 38898 39200
rect 20 856 38898 39144
rect 130 800 11554 856
rect 11722 800 23790 856
rect 23958 800 35382 856
rect 35550 800 38898 856
<< metal3 >>
rect 0 37408 800 37528
rect 39200 33328 40000 33448
rect 0 25168 800 25288
rect 39200 21088 40000 21208
rect 0 12248 800 12368
rect 39200 8168 40000 8288
<< obsm3 >>
rect 880 37328 39200 37569
rect 800 33528 39200 37328
rect 800 33248 39120 33528
rect 800 25368 39200 33248
rect 880 25088 39200 25368
rect 800 21288 39200 25088
rect 800 21008 39120 21288
rect 800 12448 39200 21008
rect 880 12168 39200 12448
rect 800 8368 39200 12168
rect 800 8088 39120 8368
rect 800 2143 39200 8088
<< metal4 >>
rect 4208 2128 4528 37584
rect 4868 2128 5188 37584
rect 34928 2128 35248 37584
rect 35588 2128 35908 37584
<< obsm4 >>
rect 34651 10915 34717 21045
<< metal5 >>
rect 1056 36642 38872 36962
rect 1056 35982 38872 36302
rect 1056 6006 38872 6326
rect 1056 5346 38872 5666
<< labels >>
rlabel metal4 s 4868 2128 5188 37584 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 35588 2128 35908 37584 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 6006 38872 6326 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 36642 38872 36962 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4208 2128 4528 37584 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 37584 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5346 38872 5666 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 35982 38872 36302 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 39200 21088 40000 21208 6 clk
port 3 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 data_in[0]
port 4 nsew signal input
rlabel metal2 s 33506 39200 33562 40000 6 data_in[1]
port 5 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 data_in[2]
port 6 nsew signal input
rlabel metal2 s 18 0 74 800 6 data_in[3]
port 7 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 data_in[4]
port 8 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 data_in[5]
port 9 nsew signal input
rlabel metal2 s 21914 39200 21970 40000 6 data_in[6]
port 10 nsew signal input
rlabel metal3 s 39200 33328 40000 33448 6 data_in[7]
port 11 nsew signal input
rlabel metal2 s 11610 0 11666 800 6 rst_n
port 12 nsew signal input
rlabel metal3 s 0 37408 800 37528 6 tx_busy
port 13 nsew signal output
rlabel metal2 s 9678 39200 9734 40000 6 tx_out
port 14 nsew signal output
rlabel metal3 s 39200 8168 40000 8288 6 tx_start
port 15 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1119524
string GDS_FILE /openlane/designs/uart_tx/runs/RUN_2025.12.11_20.26.15/results/signoff/uart_tx.magic.gds
string GDS_START 350530
<< end >>

