magic
tech sky130A
magscale 1 2
timestamp 1765482297
<< obsli1 >>
rect 1104 2159 28888 27761
<< obsm1 >>
rect 14 2128 28888 27792
<< metal2 >>
rect 7102 29200 7158 30000
rect 16118 29200 16174 30000
rect 25134 29200 25190 30000
rect 18 0 74 800
rect 9034 0 9090 800
rect 18050 0 18106 800
rect 27066 0 27122 800
<< obsm2 >>
rect 20 29144 7046 29322
rect 7214 29144 16062 29322
rect 16230 29144 25078 29322
rect 25246 29144 28594 29322
rect 20 856 28594 29144
rect 130 800 8978 856
rect 9146 800 17994 856
rect 18162 800 27010 856
rect 27178 800 28594 856
<< metal3 >>
rect 0 27888 800 28008
rect 29200 25168 30000 25288
rect 0 18368 800 18488
rect 29200 15648 30000 15768
rect 0 8848 800 8968
rect 29200 6128 30000 6248
<< obsm3 >>
rect 880 27808 29200 27978
rect 798 25368 29200 27808
rect 798 25088 29120 25368
rect 798 18568 29200 25088
rect 880 18288 29200 18568
rect 798 15848 29200 18288
rect 798 15568 29120 15848
rect 798 9048 29200 15568
rect 880 8768 29200 9048
rect 798 6328 29200 8768
rect 798 6048 29120 6328
rect 798 2143 29200 6048
<< metal4 >>
rect 4417 2128 4737 27792
rect 5077 2128 5397 27792
rect 11363 2128 11683 27792
rect 12023 2128 12343 27792
rect 18309 2128 18629 27792
rect 18969 2128 19289 27792
rect 25255 2128 25575 27792
rect 25915 2128 26235 27792
<< obsm4 >>
rect 24899 8195 24965 15741
<< metal5 >>
rect 1056 25048 28936 25368
rect 1056 24388 28936 24708
rect 1056 18656 28936 18976
rect 1056 17996 28936 18316
rect 1056 12264 28936 12584
rect 1056 11604 28936 11924
rect 1056 5872 28936 6192
rect 1056 5212 28936 5532
<< labels >>
rlabel metal4 s 5077 2128 5397 27792 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 12023 2128 12343 27792 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 18969 2128 19289 27792 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 25915 2128 26235 27792 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 5872 28936 6192 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 12264 28936 12584 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 18656 28936 18976 6 VGND
port 1 nsew ground bidirectional
rlabel metal5 s 1056 25048 28936 25368 6 VGND
port 1 nsew ground bidirectional
rlabel metal4 s 4417 2128 4737 27792 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 11363 2128 11683 27792 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 18309 2128 18629 27792 6 VPWR
port 2 nsew power bidirectional
rlabel metal4 s 25255 2128 25575 27792 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 5212 28936 5532 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 11604 28936 11924 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 17996 28936 18316 6 VPWR
port 2 nsew power bidirectional
rlabel metal5 s 1056 24388 28936 24708 6 VPWR
port 2 nsew power bidirectional
rlabel metal3 s 29200 15648 30000 15768 6 clk
port 3 nsew signal input
rlabel metal2 s 18050 0 18106 800 6 data_in[0]
port 4 nsew signal input
rlabel metal2 s 25134 29200 25190 30000 6 data_in[1]
port 5 nsew signal input
rlabel metal3 s 0 18368 800 18488 6 data_in[2]
port 6 nsew signal input
rlabel metal2 s 18 0 74 800 6 data_in[3]
port 7 nsew signal input
rlabel metal2 s 27066 0 27122 800 6 data_in[4]
port 8 nsew signal input
rlabel metal3 s 0 8848 800 8968 6 data_in[5]
port 9 nsew signal input
rlabel metal2 s 16118 29200 16174 30000 6 data_in[6]
port 10 nsew signal input
rlabel metal3 s 29200 25168 30000 25288 6 data_in[7]
port 11 nsew signal input
rlabel metal2 s 9034 0 9090 800 6 rst_n
port 12 nsew signal input
rlabel metal3 s 0 27888 800 28008 6 tx_busy
port 13 nsew signal output
rlabel metal2 s 7102 29200 7158 30000 6 tx_out
port 14 nsew signal output
rlabel metal3 s 29200 6128 30000 6248 6 tx_start
port 15 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 30000 30000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 1041146
string GDS_FILE /openlane/designs/uart_tx/runs/RUN_2025.12.11_19.43.52/results/signoff/uart_tx.magic.gds
string GDS_START 345926
<< end >>

